VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  MACRO write_qor_data STRING ;
  MACRO previous_effective_target_usage REAL ;
  MACRO achieved_target_routing_density REAL ;
  MACRO expanded_util REAL ;
END PROPERTYDEFINITIONS

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.135 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.1 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.1 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.1 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.1 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.1 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 ;
  WIDTH 0.4 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.4 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.8 ;
  WIDTH 0.4 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.4 WRONGDIRECTION ;" ;
END M8

LAYER RV
  TYPE CUT ;
END RV

LAYER AP
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END AP

LAYER M1_TEXT
  TYPE MASTERSLICE ;
END M1_TEXT

LAYER M2_TEXT
  TYPE MASTERSLICE ;
END M2_TEXT

LAYER M3_TEXT
  TYPE MASTERSLICE ;
END M3_TEXT

LAYER M4_TEXT
  TYPE MASTERSLICE ;
END M4_TEXT

LAYER M5_TEXT
  TYPE MASTERSLICE ;
END M5_TEXT

LAYER M6_TEXT
  TYPE MASTERSLICE ;
END M6_TEXT

LAYER M7_TEXT
  TYPE MASTERSLICE ;
END M7_TEXT

LAYER M8_TEXT
  TYPE MASTERSLICE ;
END M8_TEXT

LAYER VTL_N
  TYPE MASTERSLICE ;
END VTL_N

LAYER VTL_P
  TYPE MASTERSLICE ;
END VTL_P

LAYER VTH_N
  TYPE MASTERSLICE ;
END VTH_N

LAYER VTH_P
  TYPE MASTERSLICE ;
END VTH_P

LAYER VTUL_N
  TYPE MASTERSLICE ;
END VTUL_N

LAYER VTUL_P
  TYPE MASTERSLICE ;
END VTUL_P

LAYER UHVT_N
  TYPE MASTERSLICE ;
END UHVT_N

LAYER UHVT_P
  TYPE MASTERSLICE ;
END UHVT_P

LAYER PR
  TYPE MASTERSLICE ;
END PR

LAYER DIODEMY
  TYPE MASTERSLICE ;
END DIODEMY

LAYER TAP_MARKER
  TYPE MASTERSLICE ;
END TAP_MARKER

LAYER PM
  TYPE MASTERSLICE ;
END PM

LAYER PW
  TYPE MASTERSLICE ;
END PW

LAYER OD
  TYPE MASTERSLICE ;
END OD

LAYER NP
  TYPE MASTERSLICE ;
END NP

LAYER PP
  TYPE MASTERSLICE ;
END PP

LAYER NW
  TYPE MASTERSLICE ;
END NW

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE MASTERSLICE ;
END CO

LAYER GB1_5
  TYPE MASTERSLICE ;
END GB1_5

LAYER OD_18
  TYPE MASTERSLICE ;
END OD_18

LAYER OD_25
  TYPE MASTERSLICE ;
END OD_25

LAYER RPO
  TYPE MASTERSLICE ;
END RPO

LAYER RODMY
  TYPE MASTERSLICE ;
END RODMY

LAYER SRM
  TYPE MASTERSLICE ;
END SRM

LAYER CB
  TYPE MASTERSLICE ;
END CB

LAYER CB2_FC
  TYPE MASTERSLICE ;
END CB2_FC

LAYER PSUB2
  TYPE MASTERSLICE ;
END PSUB2

LAYER SR_ESD
  TYPE MASTERSLICE ;
END SR_ESD

LAYER SDI
  TYPE MASTERSLICE ;
END SDI

LAYER AP_PIN
  TYPE MASTERSLICE ;
END AP_PIN

LAYER VAR
  TYPE MASTERSLICE ;
END VAR

LAYER PO_PIN
  TYPE MASTERSLICE ;
END PO_PIN

LAYER WBDMY
  TYPE MASTERSLICE ;
END WBDMY

LAYER SRAMDMY
  TYPE MASTERSLICE ;
END SRAMDMY

LAYER ESDIMP
  TYPE MASTERSLICE ;
END ESDIMP

LAYER LVSDMY
  TYPE MASTERSLICE ;
END LVSDMY

LAYER VDDDMY
  TYPE MASTERSLICE ;
END VDDDMY

LAYER IP_BASE0
  TYPE MASTERSLICE ;
END IP_BASE0

LAYER AP_TEXT_BASE0
  TYPE MASTERSLICE ;
END AP_TEXT_BASE0

LAYER RPDMY_BASE0
  TYPE MASTERSLICE ;
END RPDMY_BASE0

LAYER RPDMY_DG1_BASE0
  TYPE MASTERSLICE ;
END RPDMY_DG1_BASE0

LAYER RH_BASE0
  TYPE MASTERSLICE ;
END RH_BASE0

LAYER DMEXCL_DUMMY1_BASE0
  TYPE MASTERSLICE ;
END DMEXCL_DUMMY1_BASE0

VIA VIA1_0_30_0_30_VH_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_0_30_0_30_VH_VX

VIA VIA1_0_30_20_20_VX_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.045 -0.045 0.045 0.045 ;
END VIA1_0_30_20_20_VX_VX

VIA VIA1_20_20_0_30_XH_VX
  LAYER M1 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_20_20_0_30_XH_VX

VIA VIA1_20_20_20_20_XX_VX
  LAYER M1 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.045 -0.045 0.045 0.045 ;
END VIA1_20_20_20_20_XX_VX

VIA VIA1_0_30_0_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_0_30_0_30_HH_VX

VIA VIA1_0_30_0_30_VV_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_0_30_0_30_VV_VX

VIA VIA1_0_30_0_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_0_30_0_30_HV_VX

VIA VIA1_0_30_5_30_VH_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_0_30_5_30_VH_VX

VIA VIA1_0_30_5_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_0_30_5_30_HH_VX

VIA VIA1_0_30_5_30_VV_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_0_30_5_30_VV_VX

VIA VIA1_0_30_5_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_0_30_5_30_HV_VX

VIA VIA1_0_30_15_30_VH_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_0_30_15_30_VH_VX

VIA VIA1_0_30_15_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_0_30_15_30_HH_VX

VIA VIA1_0_30_15_30_VV_VX
  LAYER M1 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_0_30_15_30_VV_VX

VIA VIA1_0_30_15_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_0_30_15_30_HV_VX

VIA VIA1_0_40_0_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA1_0_40_0_40_VXRECT_H

VIA VIA1_0_40_0_40_VXRECT_V
  LAYER M1 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA1_0_40_0_40_VXRECT_V

VIA VIA1_0_40_5_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA1_0_40_5_40_VXRECT_H

VIA VIA1_0_40_5_40_VXRECT_V
  LAYER M1 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA1_0_40_5_40_VXRECT_V

VIA VIA1_0_40_15_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA1_0_40_15_40_VXRECT_H

VIA VIA1_0_40_15_40_VXRECT_V
  LAYER M1 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA1_0_40_15_40_VXRECT_V

VIA VIA1_5_30_0_30_VH_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_5_30_0_30_VH_VX

VIA VIA1_5_30_0_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_5_30_0_30_HH_VX

VIA VIA1_5_30_0_30_VV_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_5_30_0_30_VV_VX

VIA VIA1_5_30_0_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_5_30_0_30_HV_VX

VIA VIA1_5_30_5_30_VH_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_5_30_5_30_VH_VX

VIA VIA1_5_30_5_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_5_30_5_30_HH_VX

VIA VIA1_5_30_5_30_VV_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_5_30_5_30_VV_VX

VIA VIA1_5_30_5_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_5_30_5_30_HV_VX

VIA VIA1_5_30_15_30_VH_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_5_30_15_30_VH_VX

VIA VIA1_5_30_15_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_5_30_15_30_HH_VX

VIA VIA1_5_30_15_30_VV_VX
  LAYER M1 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_5_30_15_30_VV_VX

VIA VIA1_5_30_15_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_5_30_15_30_HV_VX

VIA VIA1_5_40_0_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA1_5_40_0_40_VXRECT_H

VIA VIA1_5_40_0_40_VXRECT_V
  LAYER M1 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA1_5_40_0_40_VXRECT_V

VIA VIA1_5_40_5_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA1_5_40_5_40_VXRECT_H

VIA VIA1_5_40_5_40_VXRECT_V
  LAYER M1 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA1_5_40_5_40_VXRECT_V

VIA VIA1_5_40_15_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA1_5_40_15_40_VXRECT_H

VIA VIA1_5_40_15_40_VXRECT_V
  LAYER M1 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA1_5_40_15_40_VXRECT_V

VIA VIA1_15_30_0_30_VH_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_15_30_0_30_VH_VX

VIA VIA1_15_30_0_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA1_15_30_0_30_HH_VX

VIA VIA1_15_30_0_30_VV_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_15_30_0_30_VV_VX

VIA VIA1_15_30_0_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA1_15_30_0_30_HV_VX

VIA VIA1_15_30_5_30_VH_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_15_30_5_30_VH_VX

VIA VIA1_15_30_5_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA1_15_30_5_30_HH_VX

VIA VIA1_15_30_5_30_VV_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_15_30_5_30_VV_VX

VIA VIA1_15_30_5_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA1_15_30_5_30_HV_VX

VIA VIA1_15_30_15_30_VH_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_15_30_15_30_VH_VX

VIA VIA1_15_30_15_30_HH_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA1_15_30_15_30_HH_VX

VIA VIA1_15_30_15_30_VV_VX
  LAYER M1 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_15_30_15_30_VV_VX

VIA VIA1_15_30_15_30_HV_VX
  LAYER M1 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA1_15_30_15_30_HV_VX

VIA VIA1_15_40_0_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA1_15_40_0_40_VXRECT_H

VIA VIA1_15_40_0_40_VXRECT_V
  LAYER M1 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA1_15_40_0_40_VXRECT_V

VIA VIA1_15_40_5_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA1_15_40_5_40_VXRECT_H

VIA VIA1_15_40_5_40_VXRECT_V
  LAYER M1 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA1_15_40_5_40_VXRECT_V

VIA VIA1_15_40_15_40_VXRECT_H
  LAYER M1 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA1 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA1_15_40_15_40_VXRECT_H

VIA VIA1_15_40_15_40_VXRECT_V
  LAYER M1 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA1 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA1_15_40_15_40_VXRECT_V

VIA VIA2_0_30_0_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_0_30_0_30_HV_VX

VIA VIA2_0_30_0_30_VV_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_0_30_0_30_VV_VX

VIA VIA2_0_30_0_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_0_30_0_30_HH_VX

VIA VIA2_0_30_0_30_VH_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_0_30_0_30_VH_VX

VIA VIA2_0_30_5_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_0_30_5_30_HV_VX

VIA VIA2_0_30_5_30_VV_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_0_30_5_30_VV_VX

VIA VIA2_0_30_5_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_0_30_5_30_HH_VX

VIA VIA2_0_30_5_30_VH_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_0_30_5_30_VH_VX

VIA VIA2_0_30_15_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_0_30_15_30_HV_VX

VIA VIA2_0_30_15_30_VV_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_0_30_15_30_VV_VX

VIA VIA2_0_30_15_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_0_30_15_30_HH_VX

VIA VIA2_0_30_15_30_VH_VX
  LAYER M2 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_0_30_15_30_VH_VX

VIA VIA2_30_10_30_10_VXRECT_H
  LAYER M2 ;
    RECT -0.075 -0.055 0.075 0.055 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.075 -0.055 0.075 0.055 ;
END VIA2_30_10_30_10_VXRECT_H

VIA VIA2_30_10_30_10_VXRECT_V
  LAYER M2 ;
    RECT -0.055 -0.075 0.055 0.075 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.055 -0.075 0.055 0.075 ;
END VIA2_30_10_30_10_VXRECT_V

VIA VIA2_0_40_0_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA2_0_40_0_40_VXRECT_H

VIA VIA2_0_40_0_40_VXRECT_V
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA2_0_40_0_40_VXRECT_V

VIA VIA2_0_40_5_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA2_0_40_5_40_VXRECT_H

VIA VIA2_0_40_5_40_VXRECT_V
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA2_0_40_5_40_VXRECT_V

VIA VIA2_0_40_15_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA2_0_40_15_40_VXRECT_H

VIA VIA2_0_40_15_40_VXRECT_V
  LAYER M2 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA2_0_40_15_40_VXRECT_V

VIA VIA2_5_30_0_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_5_30_0_30_HV_VX

VIA VIA2_5_30_0_30_VV_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_5_30_0_30_VV_VX

VIA VIA2_5_30_0_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_5_30_0_30_HH_VX

VIA VIA2_5_30_0_30_VH_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_5_30_0_30_VH_VX

VIA VIA2_5_30_5_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_5_30_5_30_HV_VX

VIA VIA2_5_30_5_30_VV_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_5_30_5_30_VV_VX

VIA VIA2_5_30_5_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_5_30_5_30_HH_VX

VIA VIA2_5_30_5_30_VH_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_5_30_5_30_VH_VX

VIA VIA2_5_30_15_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_5_30_15_30_HV_VX

VIA VIA2_5_30_15_30_VV_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_5_30_15_30_VV_VX

VIA VIA2_5_30_15_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_5_30_15_30_HH_VX

VIA VIA2_5_30_15_30_VH_VX
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_5_30_15_30_VH_VX

VIA VIA2_5_40_0_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA2_5_40_0_40_VXRECT_H

VIA VIA2_5_40_0_40_VXRECT_V
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA2_5_40_0_40_VXRECT_V

VIA VIA2_5_40_5_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA2_5_40_5_40_VXRECT_H

VIA VIA2_5_40_5_40_VXRECT_V
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA2_5_40_5_40_VXRECT_V

VIA VIA2_5_40_15_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA2_5_40_15_40_VXRECT_H

VIA VIA2_5_40_15_40_VXRECT_V
  LAYER M2 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA2_5_40_15_40_VXRECT_V

VIA VIA2_15_30_0_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_15_30_0_30_HV_VX

VIA VIA2_15_30_0_30_VV_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA2_15_30_0_30_VV_VX

VIA VIA2_15_30_0_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_15_30_0_30_HH_VX

VIA VIA2_15_30_0_30_VH_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA2_15_30_0_30_VH_VX

VIA VIA2_15_30_5_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_15_30_5_30_HV_VX

VIA VIA2_15_30_5_30_VV_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA2_15_30_5_30_VV_VX

VIA VIA2_15_30_5_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_15_30_5_30_HH_VX

VIA VIA2_15_30_5_30_VH_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA2_15_30_5_30_VH_VX

VIA VIA2_15_30_15_30_HV_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_15_30_15_30_HV_VX

VIA VIA2_15_30_15_30_VV_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA2_15_30_15_30_VV_VX

VIA VIA2_15_30_15_30_HH_VX
  LAYER M2 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_15_30_15_30_HH_VX

VIA VIA2_15_30_15_30_VH_VX
  LAYER M2 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA2_15_30_15_30_VH_VX

VIA VIA2_15_40_0_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA2_15_40_0_40_VXRECT_H

VIA VIA2_15_40_0_40_VXRECT_V
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA2_15_40_0_40_VXRECT_V

VIA VIA2_15_40_5_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA2_15_40_5_40_VXRECT_H

VIA VIA2_15_40_5_40_VXRECT_V
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA2_15_40_5_40_VXRECT_V

VIA VIA2_15_40_15_40_VXRECT_H
  LAYER M2 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA2 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA2_15_40_15_40_VXRECT_H

VIA VIA2_15_40_15_40_VXRECT_V
  LAYER M2 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA2 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA2_15_40_15_40_VXRECT_V

VIA VIA3_0_30_0_30_VH_VX
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_0_30_0_30_VH_VX

VIA VIA3_0_30_0_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_0_30_0_30_HH_VX

VIA VIA3_0_30_5_30_VH_VX
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_0_30_5_30_VH_VX

VIA VIA3_0_30_5_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_0_30_5_30_HH_VX

VIA VIA3_0_30_15_30_VH_VX
  LAYER M3 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_0_30_15_30_VH_VX

VIA VIA3_0_30_15_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_0_30_15_30_HH_VX

VIA VIA3_0_40_0_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA3_0_40_0_40_VXRECT_H

VIA VIA3_0_40_0_40_VXRECT_V
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA3_0_40_0_40_VXRECT_V

VIA VIA3_30_10_30_10_VXRECT_H
  LAYER M3 ;
    RECT -0.075 -0.055 0.075 0.055 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.075 -0.055 0.075 0.055 ;
END VIA3_30_10_30_10_VXRECT_H

VIA VIA3_30_10_30_10_VXRECT_V
  LAYER M3 ;
    RECT -0.055 -0.075 0.055 0.075 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.055 -0.075 0.055 0.075 ;
END VIA3_30_10_30_10_VXRECT_V

VIA VIA3_0_40_5_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA3_0_40_5_40_VXRECT_H

VIA VIA3_0_40_5_40_VXRECT_V
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA3_0_40_5_40_VXRECT_V

VIA VIA3_0_40_15_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA3_0_40_15_40_VXRECT_H

VIA VIA3_0_40_15_40_VXRECT_V
  LAYER M3 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA3_0_40_15_40_VXRECT_V

VIA VIA3_5_30_0_30_VH_VX
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_5_30_0_30_VH_VX

VIA VIA3_5_30_0_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_5_30_0_30_HH_VX

VIA VIA3_5_30_5_30_VH_VX
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_5_30_5_30_VH_VX

VIA VIA3_5_30_5_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_5_30_5_30_HH_VX

VIA VIA3_5_30_15_30_VH_VX
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_5_30_15_30_VH_VX

VIA VIA3_5_30_15_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_5_30_15_30_HH_VX

VIA VIA3_5_40_0_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA3_5_40_0_40_VXRECT_H

VIA VIA3_5_40_0_40_VXRECT_V
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA3_5_40_0_40_VXRECT_V

VIA VIA3_5_40_5_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA3_5_40_5_40_VXRECT_H

VIA VIA3_5_40_5_40_VXRECT_V
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA3_5_40_5_40_VXRECT_V

VIA VIA3_5_40_15_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA3_5_40_15_40_VXRECT_H

VIA VIA3_5_40_15_40_VXRECT_V
  LAYER M3 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA3_5_40_15_40_VXRECT_V

VIA VIA3_15_30_0_30_VH_VX
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_15_30_0_30_VH_VX

VIA VIA3_15_30_0_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA3_15_30_0_30_HH_VX

VIA VIA3_15_30_5_30_VH_VX
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_15_30_5_30_VH_VX

VIA VIA3_15_30_5_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA3_15_30_5_30_HH_VX

VIA VIA3_15_30_15_30_VH_VX
  LAYER M3 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_15_30_15_30_VH_VX

VIA VIA3_15_30_15_30_HH_VX
  LAYER M3 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA3_15_30_15_30_HH_VX

VIA VIA3_15_40_0_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA3_15_40_0_40_VXRECT_H

VIA VIA3_15_40_0_40_VXRECT_V
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA3_15_40_0_40_VXRECT_V

VIA VIA3_15_40_5_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA3_15_40_5_40_VXRECT_H

VIA VIA3_15_40_5_40_VXRECT_V
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA3_15_40_5_40_VXRECT_V

VIA VIA3_15_40_15_40_VXRECT_H
  LAYER M3 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA3 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA3_15_40_15_40_VXRECT_H

VIA VIA3_15_40_15_40_VXRECT_V
  LAYER M3 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA3 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M4 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA3_15_40_15_40_VXRECT_V

VIA VIA4_0_30_0_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA4_0_30_0_30_HV_VX

VIA VIA4_0_30_5_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA4_0_30_5_30_HV_VX

VIA VIA4_0_30_15_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.025 0.055 0.025 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA4_0_30_15_30_HV_VX

VIA VIA4_0_40_0_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA4_0_40_0_40_VXRECT_H

VIA VIA4_0_40_0_40_VXRECT_V
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA4_0_40_0_40_VXRECT_V

VIA VIA4_0_40_5_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA4_0_40_5_40_VXRECT_H

VIA VIA4_30_10_30_10_VXRECT_H
  LAYER M4 ;
    RECT -0.075 -0.055 0.075 0.055 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.075 -0.055 0.075 0.055 ;
END VIA4_30_10_30_10_VXRECT_H

VIA VIA4_30_10_30_10_VXRECT_V
  LAYER M4 ;
    RECT -0.055 -0.075 0.055 0.075 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.055 -0.075 0.055 0.075 ;
END VIA4_30_10_30_10_VXRECT_V

VIA VIA4_0_40_5_40_VXRECT_V
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA4_0_40_5_40_VXRECT_V

VIA VIA4_0_40_15_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA4_0_40_15_40_VXRECT_H

VIA VIA4_0_40_15_40_VXRECT_V
  LAYER M4 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA4_0_40_15_40_VXRECT_V

VIA VIA4_5_30_0_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA4_5_30_0_30_HV_VX

VIA VIA4_5_30_5_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA4_5_30_5_30_HV_VX

VIA VIA4_5_30_15_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA4_5_30_15_30_HV_VX

VIA VIA4_5_40_0_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA4_5_40_0_40_VXRECT_H

VIA VIA4_5_40_0_40_VXRECT_V
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA4_5_40_0_40_VXRECT_V

VIA VIA4_5_40_5_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA4_5_40_5_40_VXRECT_H

VIA VIA4_5_40_5_40_VXRECT_V
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA4_5_40_5_40_VXRECT_V

VIA VIA4_5_40_15_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA4_5_40_15_40_VXRECT_H

VIA VIA4_5_40_15_40_VXRECT_V
  LAYER M4 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA4_5_40_15_40_VXRECT_V

VIA VIA4_15_30_0_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
END VIA4_15_30_0_30_HV_VX

VIA VIA4_15_30_5_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA4_15_30_5_30_HV_VX

VIA VIA4_15_30_15_30_HV_VX
  LAYER M4 ;
    RECT -0.055 -0.04 0.055 0.04 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
END VIA4_15_30_15_30_HV_VX

VIA VIA4_15_40_0_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA4_15_40_0_40_VXRECT_H

VIA VIA4_15_40_0_40_VXRECT_V
  LAYER M4 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA4_15_40_0_40_VXRECT_V

VIA VIA4_15_40_5_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA4_15_40_5_40_VXRECT_H

VIA VIA4_15_40_15_40_VXRECT_H
  LAYER M4 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA4 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA4_15_40_15_40_VXRECT_H

VIA VIA4_15_40_15_40_VXRECT_V
  LAYER M4 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA4 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA4_15_40_15_40_VXRECT_V

VIA VIA5_0_30_0_30_VH_VX
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA5_0_30_0_30_VH_VX

VIA VIA5_0_30_5_30_VH_VX
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA5_0_30_5_30_VH_VX

VIA VIA5_0_30_15_30_VH_VX
  LAYER M5 ;
    RECT -0.025 -0.055 0.025 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA5_0_30_15_30_VH_VX

VIA VIA5_30_10_30_10_VXRECT_H
  LAYER M5 ;
    RECT -0.075 -0.055 0.075 0.055 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.075 -0.055 0.075 0.055 ;
END VIA5_30_10_30_10_VXRECT_H

VIA VIA5_30_10_30_10_VXRECT_V
  LAYER M5 ;
    RECT -0.055 -0.075 0.055 0.075 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.055 -0.075 0.055 0.075 ;
END VIA5_30_10_30_10_VXRECT_V

VIA VIA5_0_40_0_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA5_0_40_0_40_VXRECT_H

VIA VIA5_0_40_0_40_VXRECT_V
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA5_0_40_0_40_VXRECT_V

VIA VIA5_0_40_5_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA5_0_40_5_40_VXRECT_H

VIA VIA5_0_40_5_40_VXRECT_V
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA5_0_40_5_40_VXRECT_V

VIA VIA5_0_40_15_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.025 0.105 0.025 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA5_0_40_15_40_VXRECT_H

VIA VIA5_0_40_15_40_VXRECT_V
  LAYER M5 ;
    RECT -0.025 -0.105 0.025 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA5_0_40_15_40_VXRECT_V

VIA VIA5_5_30_0_30_VH_VX
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA5_5_30_0_30_VH_VX

VIA VIA5_5_30_5_30_VH_VX
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA5_5_30_5_30_VH_VX

VIA VIA5_5_30_15_30_VH_VX
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA5_5_30_15_30_VH_VX

VIA VIA5_5_40_0_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA5_5_40_0_40_VXRECT_H

VIA VIA5_5_40_0_40_VXRECT_V
  LAYER M5 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA5_5_40_0_40_VXRECT_V

VIA VIA5_5_40_5_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA5_5_40_5_40_VXRECT_H

VIA VIA5_5_40_5_40_VXRECT_V
  LAYER M5 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA5_5_40_5_40_VXRECT_V

VIA VIA5_5_40_15_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.03 0.105 0.03 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA5_5_40_15_40_VXRECT_H

VIA VIA5_5_40_15_40_VXRECT_V
  LAYER M5 ;
    RECT -0.03 -0.105 0.03 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA5_5_40_15_40_VXRECT_V

VIA VIA5_15_30_0_30_VH_VX
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.025 0.055 0.025 ;
END VIA5_15_30_0_30_VH_VX

VIA VIA5_15_30_5_30_VH_VX
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA5_15_30_5_30_VH_VX

VIA VIA5_15_30_15_30_VH_VX
  LAYER M5 ;
    RECT -0.04 -0.055 0.04 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.04 0.055 0.04 ;
END VIA5_15_30_15_30_VH_VX

VIA VIA5_15_40_0_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.025 0.105 0.025 ;
END VIA5_15_40_0_40_VXRECT_H

VIA VIA5_15_40_0_40_VXRECT_V
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.025 -0.105 0.025 0.105 ;
END VIA5_15_40_0_40_VXRECT_V

VIA VIA5_15_40_5_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.03 0.105 0.03 ;
END VIA5_15_40_5_40_VXRECT_H

VIA VIA5_15_40_5_40_VXRECT_V
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.03 -0.105 0.03 0.105 ;
END VIA5_15_40_5_40_VXRECT_V

VIA VIA5_15_40_15_40_VXRECT_H
  LAYER M5 ;
    RECT -0.105 -0.04 0.105 0.04 ;
  LAYER VIA5 ;
    RECT -0.065 -0.025 0.065 0.025 ;
  LAYER M6 ;
    RECT -0.105 -0.04 0.105 0.04 ;
END VIA5_15_40_15_40_VXRECT_H

VIA VIA5_15_40_15_40_VXRECT_V
  LAYER M5 ;
    RECT -0.04 -0.105 0.04 0.105 ;
  LAYER VIA5 ;
    RECT -0.025 -0.065 0.025 0.065 ;
  LAYER M6 ;
    RECT -0.04 -0.105 0.04 0.105 ;
END VIA5_15_40_15_40_VXRECT_V

VIA VIA6_20_80_20_80_HV_VZ_F0
  LAYER M6 ;
    RECT -0.26 -0.2 0.26 0.2 ;
  LAYER VIA6 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M7 ;
    RECT -0.2 -0.26 0.2 0.26 ;
END VIA6_20_80_20_80_HV_VZ_F0

VIA VIA6_20_80_20_80_HV_VZ_F0_fat
  LAYER M6 ;
    RECT -0.26 -0.2 0.26 0.2 ;
  LAYER VIA6 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M7 ;
    RECT -0.26 -0.2 0.26 0.2 ;
END VIA6_20_80_20_80_HV_VZ_F0_fat

VIA VIA7_20_80_20_80_VH_VZ_F0
  LAYER M7 ;
    RECT -0.2 -0.26 0.2 0.26 ;
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.26 -0.2 0.26 0.2 ;
END VIA7_20_80_20_80_VH_VZ_F0

VIA VIA7_20_80_20_80_VH_VZ_F0_fat
  LAYER M7 ;
    RECT -0.26 -0.2 0.26 0.2 ;
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.26 -0.2 0.26 0.2 ;
END VIA7_20_80_20_80_VH_VZ_F0_fat

VIA RV_500_500_500_500_XX
  LAYER M8 ;
    RECT -2 -2 2 2 ;
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER AP ;
    RECT -2 -2 2 2 ;
END RV_500_500_500_500_XX

SITE sc12mc_cln28hpm
  CLASS CORE ;
  SIZE 0.135 BY 1.2 ;
END sc12mc_cln28hpm

MACRO DFFRPQL_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN DFFRPQL_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.165 0.295 0.235 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0105 ;
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.525 0.705 2.525 0.495 2.555 0.495 2.555 0.425 2.44 0.425 2.44 0.495 2.465 0.495 2.465 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0084 ;
  END CK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.985 0.625 1.035 0.675 ;
        RECT 1.82 0.625 1.95 0.675 ;
      LAYER M1 ;
        POLYGON 1.99 0.685 1.99 0.615 1.86 0.615 1.86 0.525 1.78 0.525 1.78 0.685 ;
        RECT 0.975 0.465 1.045 0.74 ;
      LAYER M2 ;
        RECT 0.935 0.625 2 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0077 LAYER M1 ;
    ANTENNAGATEAREA 0.0224 LAYER M2 ;
    ANTENNAGATEAREA 0.0224 LAYER M3 ;
    ANTENNAGATEAREA 0.0224 LAYER M4 ;
    ANTENNAGATEAREA 0.0224 LAYER M5 ;
    ANTENNAGATEAREA 0.0224 LAYER M6 ;
    ANTENNAGATEAREA 0.0224 LAYER M7 ;
    ANTENNAGATEAREA 0.0224 LAYER M8 ;
    ANTENNAGATEAREA 0.0224 LAYER AP ;
    ANTENNAMAXAREACAR 2.844156 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.8441558 LAYER VIA1 ;
  END R
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.32 0.945 2.32 0.805 2.39 0.805 2.39 0.375 2.32 0.375 2.32 0.235 2.27 0.235 2.27 0.425 2.335 0.425 2.335 0.755 2.27 0.755 2.27 0.945 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
      LAYER M1 ;
        POLYGON 2.835 1.235 2.835 1.165 2.61 1.165 2.61 0.925 2.54 0.925 2.54 1.165 2.195 1.165 2.195 0.88 2.125 0.88 2.125 1.165 1.925 1.165 1.925 0.905 1.855 0.905 1.855 1.165 0.845 1.165 0.845 0.775 0.775 0.775 0.775 1.165 0.17 1.165 0.17 0.79 0.1 0.79 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.835 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.285 1.79 0.035 2.125 0.035 2.125 0.255 2.195 0.255 2.195 0.035 2.53 0.035 2.53 0.165 2.6 0.165 2.6 0.035 2.835 0.035 2.835 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.19 0.17 0.19 0.17 0.035 0.775 0.035 0.775 0.18 0.845 0.18 0.845 0.035 1.045 0.035 1.045 0.19 1.115 0.19 1.115 0.035 1.72 0.035 1.72 0.285 ;
      LAYER M2 ;
        RECT 0 -0.065 2.835 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.615 1.105 1.615 0.975 1.785 0.975 1.785 0.925 1.565 0.925 1.565 1.055 1.36 1.055 1.36 1.105 ;
      POLYGON 0.375 1.105 0.375 0.975 0.675 0.975 0.675 0.925 0.305 0.925 0.305 1.105 ;
      POLYGON 2.725 1.095 2.725 0.955 2.795 0.955 2.795 0.225 2.735 0.225 2.735 0.1 2.665 0.1 2.665 0.225 2.585 0.225 2.585 0.275 2.745 0.275 2.745 0.905 2.675 0.905 2.675 1.095 ;
      POLYGON 2.05 1.095 2.05 0.81 2.22 0.81 2.22 0.585 2.27 0.585 2.27 0.515 2.22 0.515 2.22 0.325 2.065 0.325 2.065 0.095 1.985 0.095 1.985 0.175 2.015 0.175 2.015 0.375 2.17 0.375 2.17 0.76 1.71 0.76 1.71 0.62 1.66 0.62 1.66 0.81 2 0.81 2 1.095 ;
      POLYGON 1.105 1.03 1.105 0.89 1.325 0.89 1.325 0.985 1.375 0.985 1.375 0.84 1.24 0.84 1.24 0.345 0.97 0.345 0.97 0.12 0.92 0.12 0.92 0.345 0.72 0.345 0.72 0.535 0.77 0.535 0.77 0.395 1.19 0.395 1.19 0.84 1.055 0.84 1.055 1.03 ;
      POLYGON 2.465 1.015 2.465 0.935 2.49 0.935 2.49 0.845 2.66 0.845 2.66 0.325 2.515 0.325 2.515 0.225 2.465 0.225 2.465 0.1 2.395 0.1 2.395 0.275 2.465 0.275 2.465 0.375 2.61 0.375 2.61 0.795 2.44 0.795 2.44 0.885 2.395 0.885 2.395 1.015 ;
      POLYGON 1.51 0.985 1.51 0.55 1.63 0.55 1.63 0.475 2.065 0.475 2.065 0.595 2.115 0.595 2.115 0.425 1.915 0.425 1.915 0.185 1.865 0.185 1.865 0.425 1.58 0.425 1.58 0.5 1.375 0.5 1.375 0.345 1.325 0.345 1.325 0.55 1.46 0.55 1.46 0.985 ;
      POLYGON 0.565 0.855 0.565 0.68 0.905 0.68 0.905 0.49 0.855 0.49 0.855 0.63 0.36 0.63 0.36 0.16 0.595 0.16 0.595 0.11 0.31 0.11 0.31 0.68 0.515 0.68 0.515 0.855 ;
      RECT 0.225 0.785 0.45 0.855 ;
      POLYGON 1.51 0.43 1.51 0.275 1.665 0.275 1.665 0.205 1.46 0.205 1.46 0.43 ;
      POLYGON 0.5 0.415 0.5 0.275 0.68 0.275 0.68 0.225 0.45 0.225 0.45 0.415 ;
      POLYGON 1.39 0.275 1.39 0.225 1.23 0.225 1.23 0.145 1.605 0.145 1.605 0.095 1.18 0.095 1.18 0.275 ;
    LAYER M2 ;
      RECT 0.445 0.925 2.505 0.975 ;
      RECT 0.45 0.225 2.795 0.275 ;
    LAYER VIA1 ;
      RECT 2.405 0.925 2.455 0.975 ;
      RECT 1.605 0.925 1.735 0.975 ;
      RECT 0.495 0.925 0.625 0.975 ;
      RECT 2.625 0.225 2.755 0.275 ;
      RECT 1.22 0.225 1.35 0.275 ;
      RECT 0.5 0.225 0.63 0.275 ;
  END
END DFFRPQL_X1M_A12TUL_C35

MACRO DFFRPQ_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN DFFRPQ_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.635 0.625 0.635 0.395 0.58 0.395 0.58 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.705 0.37 0.495 0.525 0.495 0.525 0.425 0.28 0.425 0.28 0.495 0.3 0.495 0.3 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0091 ;
  END CK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.39 0.625 1.44 0.675 ;
        RECT 2.2 0.625 2.25 0.675 ;
      LAYER M1 ;
        RECT 2.195 0.475 2.255 0.715 ;
        RECT 1.38 0.495 1.45 0.755 ;
      LAYER M2 ;
        RECT 1.34 0.625 2.3 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00805 LAYER M1 ;
    ANTENNAGATEAREA 0.035 LAYER M2 ;
    ANTENNAGATEAREA 0.035 LAYER M3 ;
    ANTENNAGATEAREA 0.035 LAYER M4 ;
    ANTENNAGATEAREA 0.035 LAYER M5 ;
    ANTENNAGATEAREA 0.035 LAYER M6 ;
    ANTENNAGATEAREA 0.035 LAYER M7 ;
    ANTENNAGATEAREA 0.035 LAYER M8 ;
    ANTENNAGATEAREA 0.035 LAYER AP ;
    ANTENNAMAXAREACAR 1.78882 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.310559 LAYER VIA1 ;
  END R
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.725 1.045 2.725 0.905 2.795 0.905 2.795 0.295 2.725 0.295 2.725 0.155 2.675 0.155 2.675 0.345 2.74 0.345 2.74 0.855 2.675 0.855 2.675 1.045 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
      LAYER M1 ;
        POLYGON 2.835 1.235 2.835 1.165 2.6 1.165 2.6 0.775 2.53 0.775 2.53 1.165 2.335 1.165 2.335 0.905 2.255 0.905 2.255 1.165 1.255 1.165 1.255 0.81 1.18 0.81 1.18 1.165 0.575 1.165 0.575 0.76 0.505 0.76 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.835 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
      LAYER M1 ;
        POLYGON 2.6 0.355 2.6 0.035 2.835 0.035 2.835 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.18 0.305 0.18 0.305 0.035 0.505 0.035 0.505 0.315 0.575 0.315 0.575 0.035 1.18 0.035 1.18 0.3 1.25 0.3 1.25 0.035 1.45 0.035 1.45 0.305 1.52 0.305 1.52 0.035 2.125 0.035 2.125 0.285 2.195 0.285 2.195 0.035 2.53 0.035 2.53 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.835 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.89 1.115 1.89 0.925 1.665 0.925 1.665 0.975 1.84 0.975 1.84 1.065 1.75 1.065 1.75 1.115 ;
      POLYGON 1.11 1.115 1.11 0.925 0.88 0.925 0.88 0.975 1.06 0.975 1.06 1.065 0.69 1.065 0.69 1.115 ;
      POLYGON 0.43 1.1 0.43 0.775 0.225 0.775 0.225 0.375 0.43 0.375 0.43 0.1 0.38 0.1 0.38 0.325 0.175 0.325 0.175 0.825 0.38 0.825 0.38 1.1 ;
      POLYGON 0.16 1.085 0.16 0.895 0.09 0.895 0.09 0.275 0.175 0.275 0.175 0.105 0.095 0.105 0.095 0.225 0.04 0.225 0.04 0.945 0.11 0.945 0.11 1.085 ;
      POLYGON 1.51 1.015 1.51 0.875 1.78 0.875 1.78 0.625 1.645 0.625 1.645 0.375 1.375 0.375 1.375 0.135 1.325 0.135 1.325 0.375 1.12 0.375 1.12 0.575 1.17 0.575 1.17 0.425 1.595 0.425 1.595 0.675 1.73 0.675 1.73 0.825 1.46 0.825 1.46 1.015 ;
      POLYGON 0.7 0.945 0.7 0.775 0.785 0.775 0.785 0.835 0.835 0.835 0.835 0.725 0.65 0.725 0.65 0.945 ;
      POLYGON 2.455 0.865 2.455 0.695 2.66 0.695 2.66 0.425 2.455 0.425 2.455 0.115 2.405 0.115 2.405 0.475 2.61 0.475 2.61 0.645 2.405 0.645 2.405 0.785 2.115 0.785 2.115 0.645 2.065 0.645 2.065 0.835 2.405 0.835 2.405 0.865 ;
      POLYGON 1.915 0.855 1.915 0.405 2.305 0.405 2.305 0.595 2.54 0.595 2.54 0.525 2.355 0.525 2.355 0.355 2.32 0.355 2.32 0.185 2.27 0.185 2.27 0.355 1.78 0.355 1.78 0.215 1.73 0.215 1.73 0.405 1.865 0.405 1.865 0.855 ;
      POLYGON 0.97 0.805 0.97 0.705 1.305 0.705 1.305 0.495 1.255 0.495 1.255 0.655 0.97 0.655 0.97 0.525 0.75 0.525 0.75 0.325 0.835 0.325 0.835 0.15 1 0.15 1 0.1 0.785 0.1 0.785 0.275 0.7 0.275 0.7 0.575 0.92 0.575 0.92 0.805 ;
      POLYGON 1.04 0.475 1.04 0.225 0.905 0.225 0.905 0.275 0.99 0.275 0.99 0.425 0.82 0.425 0.82 0.475 ;
      POLYGON 1.655 0.315 1.655 0.135 2.03 0.135 2.03 0.085 1.585 0.085 1.585 0.315 ;
      RECT 1.85 0.2 2.065 0.28 ;
    LAYER M2 ;
      RECT 0.33 0.925 1.885 0.975 ;
      RECT 0.04 0.225 1.695 0.275 ;
    LAYER VIA1 ;
      RECT 1.705 0.925 1.835 0.975 ;
      RECT 0.93 0.925 1.06 0.975 ;
      RECT 0.38 0.925 0.43 0.975 ;
      RECT 1.595 0.225 1.645 0.275 ;
      RECT 0.95 0.225 1 0.275 ;
      RECT 0.08 0.225 0.13 0.275 ;
  END
END DFFRPQ_X1M_A12TUL_C35

MACRO DFFRPQ_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN DFFRPQ_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.97 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.635 0.625 0.635 0.395 0.58 0.395 0.58 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.705 0.37 0.495 0.525 0.495 0.525 0.425 0.28 0.425 0.28 0.495 0.3 0.495 0.3 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0126 ;
  END CK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.39 0.625 1.44 0.675 ;
        RECT 2.2 0.625 2.25 0.675 ;
      LAYER M1 ;
        RECT 2.195 0.475 2.255 0.715 ;
        RECT 1.38 0.495 1.45 0.755 ;
      LAYER M2 ;
        RECT 1.34 0.625 2.3 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00805 LAYER M1 ;
    ANTENNAGATEAREA 0.035 LAYER M2 ;
    ANTENNAGATEAREA 0.035 LAYER M3 ;
    ANTENNAGATEAREA 0.035 LAYER M4 ;
    ANTENNAGATEAREA 0.035 LAYER M5 ;
    ANTENNAGATEAREA 0.035 LAYER M6 ;
    ANTENNAGATEAREA 0.035 LAYER M7 ;
    ANTENNAGATEAREA 0.035 LAYER M8 ;
    ANTENNAGATEAREA 0.035 LAYER AP ;
    ANTENNAMAXAREACAR 1.78882 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.310559 LAYER VIA1 ;
  END R
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.725 1.015 2.725 0.875 2.93 0.875 2.93 0.325 2.725 0.325 2.725 0.185 2.675 0.185 2.675 0.375 2.875 0.375 2.875 0.825 2.675 0.825 2.675 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
      LAYER M1 ;
        POLYGON 2.97 1.235 2.97 1.165 2.87 1.165 2.87 0.925 2.8 0.925 2.8 1.165 2.6 1.165 2.6 0.775 2.53 0.775 2.53 1.165 2.335 1.165 2.335 0.905 2.255 0.905 2.255 1.165 1.25 1.165 1.25 0.81 1.18 0.81 1.18 1.165 0.575 1.165 0.575 0.76 0.505 0.76 0.505 1.165 0.305 1.165 0.305 0.9 0.235 0.9 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.97 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
      LAYER M1 ;
        POLYGON 2.6 0.355 2.6 0.035 2.8 0.035 2.8 0.275 2.87 0.275 2.87 0.035 2.97 0.035 2.97 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.18 0.305 0.18 0.305 0.035 0.505 0.035 0.505 0.315 0.575 0.315 0.575 0.035 1.18 0.035 1.18 0.305 1.25 0.305 1.25 0.035 1.45 0.035 1.45 0.305 1.52 0.305 1.52 0.035 2.125 0.035 2.125 0.28 2.195 0.28 2.195 0.035 2.53 0.035 2.53 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.97 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.89 1.115 1.89 0.925 1.665 0.925 1.665 0.975 1.84 0.975 1.84 1.065 1.75 1.065 1.75 1.115 ;
      POLYGON 1.11 1.115 1.11 0.925 0.88 0.925 0.88 0.975 1.06 0.975 1.06 1.065 0.69 1.065 0.69 1.115 ;
      POLYGON 0.16 1.085 0.16 0.895 0.09 0.895 0.09 0.275 0.175 0.275 0.175 0.105 0.095 0.105 0.095 0.225 0.04 0.225 0.04 0.945 0.11 0.945 0.11 1.085 ;
      POLYGON 0.43 1.07 0.43 0.775 0.225 0.775 0.225 0.375 0.43 0.375 0.43 0.11 0.38 0.11 0.38 0.325 0.175 0.325 0.175 0.825 0.38 0.825 0.38 1.07 ;
      POLYGON 1.51 1.015 1.51 0.875 1.78 0.875 1.78 0.555 1.645 0.555 1.645 0.375 1.375 0.375 1.375 0.135 1.325 0.135 1.325 0.375 1.12 0.375 1.12 0.585 1.17 0.585 1.17 0.425 1.595 0.425 1.595 0.605 1.73 0.605 1.73 0.825 1.46 0.825 1.46 1.015 ;
      POLYGON 0.7 0.945 0.7 0.775 0.785 0.775 0.785 0.835 0.835 0.835 0.835 0.725 0.65 0.725 0.65 0.945 ;
      POLYGON 2.455 0.865 2.455 0.695 2.66 0.695 2.66 0.585 2.81 0.585 2.81 0.515 2.66 0.515 2.66 0.425 2.455 0.425 2.455 0.135 2.405 0.135 2.405 0.475 2.61 0.475 2.61 0.645 2.405 0.645 2.405 0.785 2.115 0.785 2.115 0.645 2.065 0.645 2.065 0.835 2.405 0.835 2.405 0.865 ;
      POLYGON 1.915 0.855 1.915 0.405 2.305 0.405 2.305 0.595 2.54 0.595 2.54 0.525 2.355 0.525 2.355 0.355 2.32 0.355 2.32 0.18 2.27 0.18 2.27 0.355 1.78 0.355 1.78 0.215 1.73 0.215 1.73 0.405 1.865 0.405 1.865 0.855 ;
      POLYGON 0.97 0.805 0.97 0.705 1.305 0.705 1.305 0.495 1.255 0.495 1.255 0.655 0.97 0.655 0.97 0.525 0.75 0.525 0.75 0.325 0.835 0.325 0.835 0.15 1 0.15 1 0.1 0.785 0.1 0.785 0.275 0.7 0.275 0.7 0.575 0.92 0.575 0.92 0.805 ;
      POLYGON 1.04 0.475 1.04 0.225 0.905 0.225 0.905 0.275 0.99 0.275 0.99 0.425 0.82 0.425 0.82 0.475 ;
      POLYGON 1.655 0.315 1.655 0.135 2.03 0.135 2.03 0.085 1.585 0.085 1.585 0.315 ;
      RECT 1.845 0.195 2.07 0.275 ;
    LAYER M2 ;
      RECT 0.33 0.925 1.885 0.975 ;
      RECT 0.04 0.225 1.695 0.275 ;
    LAYER VIA1 ;
      RECT 1.705 0.925 1.835 0.975 ;
      RECT 0.93 0.925 1.06 0.975 ;
      RECT 0.38 0.925 0.43 0.975 ;
      RECT 1.595 0.225 1.645 0.275 ;
      RECT 0.95 0.225 1 0.275 ;
      RECT 0.08 0.225 0.13 0.275 ;
  END
END DFFRPQ_X2M_A12TUL_C35

MACRO DFFRPQ_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN DFFRPQ_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.635 0.625 0.635 0.395 0.58 0.395 0.58 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.705 0.37 0.495 0.525 0.495 0.525 0.425 0.28 0.425 0.28 0.495 0.3 0.495 0.3 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END CK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.39 0.625 1.44 0.675 ;
        RECT 2.2 0.625 2.25 0.675 ;
      LAYER M1 ;
        RECT 2.195 0.475 2.255 0.715 ;
        RECT 1.38 0.495 1.45 0.755 ;
      LAYER M2 ;
        RECT 1.34 0.625 2.3 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00805 LAYER M1 ;
    ANTENNAGATEAREA 0.03605 LAYER M2 ;
    ANTENNAGATEAREA 0.03605 LAYER M3 ;
    ANTENNAGATEAREA 0.03605 LAYER M4 ;
    ANTENNAGATEAREA 0.03605 LAYER M5 ;
    ANTENNAGATEAREA 0.03605 LAYER M6 ;
    ANTENNAGATEAREA 0.03605 LAYER M7 ;
    ANTENNAGATEAREA 0.03605 LAYER M8 ;
    ANTENNAGATEAREA 0.03605 LAYER AP ;
    ANTENNAMAXAREACAR 1.78882 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.310559 LAYER VIA1 ;
  END R
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.86 1.015 2.86 0.875 3.08 0.875 3.08 1 3.13 1 3.13 0.875 3.335 0.875 3.335 0.325 3.13 0.325 3.13 0.2 3.08 0.2 3.08 0.325 2.86 0.325 2.86 0.185 2.81 0.185 2.81 0.375 3.28 0.375 3.28 0.825 2.81 0.825 2.81 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
      LAYER M1 ;
        POLYGON 3.375 1.235 3.375 1.165 3.275 1.165 3.275 0.925 3.205 0.925 3.205 1.165 3.005 1.165 3.005 0.925 2.935 0.925 2.935 1.165 2.735 1.165 2.735 0.775 2.665 0.775 2.665 1.165 2.465 1.165 2.465 0.905 2.395 0.905 2.395 1.165 2.335 1.165 2.335 0.905 2.255 0.905 2.255 1.165 1.25 1.165 1.25 0.81 1.18 0.81 1.18 1.165 0.575 1.165 0.575 0.76 0.505 0.76 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.375 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
      LAYER M1 ;
        POLYGON 2.735 0.355 2.735 0.035 2.935 0.035 2.935 0.275 3.005 0.275 3.005 0.035 3.205 0.035 3.205 0.275 3.275 0.275 3.275 0.035 3.375 0.035 3.375 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.26 0.305 0.26 0.305 0.035 0.505 0.035 0.505 0.31 0.575 0.31 0.575 0.035 1.18 0.035 1.18 0.305 1.25 0.305 1.25 0.035 1.45 0.035 1.45 0.305 1.52 0.305 1.52 0.035 2.125 0.035 2.125 0.28 2.195 0.28 2.195 0.035 2.395 0.035 2.395 0.285 2.465 0.285 2.465 0.035 2.665 0.035 2.665 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 3.375 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.89 1.115 1.89 0.925 1.665 0.925 1.665 0.975 1.84 0.975 1.84 1.065 1.75 1.065 1.75 1.115 ;
      POLYGON 1.11 1.115 1.11 0.925 0.88 0.925 0.88 0.975 1.06 0.975 1.06 1.065 0.69 1.065 0.69 1.115 ;
      POLYGON 0.43 1.095 0.43 0.775 0.225 0.775 0.225 0.375 0.43 0.375 0.43 0.105 0.38 0.105 0.38 0.325 0.175 0.325 0.175 0.825 0.38 0.825 0.38 1.095 ;
      POLYGON 0.16 1.085 0.16 0.895 0.09 0.895 0.09 0.275 0.175 0.275 0.175 0.115 0.095 0.115 0.095 0.225 0.04 0.225 0.04 0.945 0.11 0.945 0.11 1.085 ;
      POLYGON 1.51 1.015 1.51 0.875 1.78 0.875 1.78 0.555 1.645 0.555 1.645 0.375 1.375 0.375 1.375 0.165 1.325 0.165 1.325 0.375 1.12 0.375 1.12 0.585 1.17 0.585 1.17 0.425 1.595 0.425 1.595 0.605 1.73 0.605 1.73 0.825 1.46 0.825 1.46 1.015 ;
      POLYGON 0.7 0.945 0.7 0.775 0.785 0.775 0.785 0.835 0.835 0.835 0.835 0.725 0.65 0.725 0.65 0.945 ;
      POLYGON 2.59 0.925 2.59 0.695 2.795 0.695 2.795 0.575 3.22 0.575 3.22 0.525 2.795 0.525 2.795 0.425 2.59 0.425 2.59 0.175 2.54 0.175 2.54 0.475 2.745 0.475 2.745 0.645 2.54 0.645 2.54 0.785 2.115 0.785 2.115 0.645 2.065 0.645 2.065 0.835 2.54 0.835 2.54 0.925 ;
      POLYGON 1.915 0.855 1.915 0.405 2.405 0.405 2.405 0.595 2.675 0.595 2.675 0.525 2.455 0.525 2.455 0.355 2.32 0.355 2.32 0.18 2.27 0.18 2.27 0.355 1.78 0.355 1.78 0.215 1.73 0.215 1.73 0.405 1.865 0.405 1.865 0.855 ;
      POLYGON 0.97 0.805 0.97 0.71 1.31 0.71 1.31 0.495 1.26 0.495 1.26 0.66 0.97 0.66 0.97 0.525 0.75 0.525 0.75 0.325 0.835 0.325 0.835 0.15 1 0.15 1 0.1 0.785 0.1 0.785 0.275 0.7 0.275 0.7 0.575 0.92 0.575 0.92 0.805 ;
      POLYGON 1.04 0.475 1.04 0.225 0.905 0.225 0.905 0.275 0.99 0.275 0.99 0.425 0.82 0.425 0.82 0.475 ;
      POLYGON 1.655 0.315 1.655 0.135 2.03 0.135 2.03 0.085 1.585 0.085 1.585 0.315 ;
      RECT 1.845 0.195 2.07 0.275 ;
    LAYER M2 ;
      RECT 0.33 0.925 1.885 0.975 ;
      RECT 0.04 0.225 1.695 0.275 ;
    LAYER VIA1 ;
      RECT 1.705 0.925 1.835 0.975 ;
      RECT 0.93 0.925 1.06 0.975 ;
      RECT 0.38 0.925 0.43 0.975 ;
      RECT 1.595 0.225 1.645 0.275 ;
      RECT 0.95 0.225 1 0.275 ;
      RECT 0.08 0.225 0.13 0.275 ;
  END
END DFFRPQ_X4M_A12TUL_C35

MACRO DFFRPQ_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN DFFRPQ_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.105 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.635 0.625 0.635 0.395 0.58 0.395 0.58 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.705 0.37 0.495 0.525 0.495 0.525 0.425 0.28 0.425 0.28 0.495 0.3 0.495 0.3 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.014 ;
  END CK
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.39 0.625 1.44 0.675 ;
        RECT 2.2 0.625 2.25 0.675 ;
      LAYER M1 ;
        RECT 2.195 0.475 2.255 0.715 ;
        RECT 1.38 0.495 1.45 0.755 ;
      LAYER M2 ;
        RECT 1.34 0.625 2.305 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00805 LAYER M1 ;
    ANTENNAGATEAREA 0.03605 LAYER M2 ;
    ANTENNAGATEAREA 0.03605 LAYER M3 ;
    ANTENNAGATEAREA 0.03605 LAYER M4 ;
    ANTENNAGATEAREA 0.03605 LAYER M5 ;
    ANTENNAGATEAREA 0.03605 LAYER M6 ;
    ANTENNAGATEAREA 0.03605 LAYER M7 ;
    ANTENNAGATEAREA 0.03605 LAYER M8 ;
    ANTENNAGATEAREA 0.03605 LAYER AP ;
    ANTENNAMAXAREACAR 1.78882 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.310559 LAYER VIA1 ;
  END R
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.725 1.015 2.725 0.875 2.945 0.875 2.945 1 2.995 1 2.995 0.875 3.065 0.875 3.065 0.325 2.995 0.325 2.995 0.2 2.945 0.2 2.945 0.325 2.725 0.325 2.725 0.185 2.675 0.185 2.675 0.375 3.01 0.375 3.01 0.825 2.675 0.825 2.675 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
      LAYER M1 ;
        POLYGON 3.105 1.235 3.105 1.165 2.87 1.165 2.87 0.925 2.8 0.925 2.8 1.165 2.6 1.165 2.6 0.775 2.53 0.775 2.53 1.165 2.335 1.165 2.335 0.905 2.255 0.905 2.255 1.165 1.25 1.165 1.25 0.81 1.18 0.81 1.18 1.165 0.575 1.165 0.575 0.76 0.505 0.76 0.505 1.165 0.305 1.165 0.305 0.9 0.235 0.9 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.105 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
      LAYER M1 ;
        POLYGON 2.6 0.355 2.6 0.035 2.8 0.035 2.8 0.275 2.87 0.275 2.87 0.035 3.105 0.035 3.105 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.26 0.305 0.26 0.305 0.035 0.505 0.035 0.505 0.315 0.575 0.315 0.575 0.035 1.18 0.035 1.18 0.305 1.25 0.305 1.25 0.035 1.45 0.035 1.45 0.305 1.52 0.305 1.52 0.035 2.125 0.035 2.125 0.28 2.195 0.28 2.195 0.035 2.53 0.035 2.53 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 3.105 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.89 1.115 1.89 0.925 1.665 0.925 1.665 0.975 1.84 0.975 1.84 1.065 1.75 1.065 1.75 1.115 ;
      POLYGON 1.11 1.115 1.11 0.925 0.88 0.925 0.88 0.975 1.06 0.975 1.06 1.065 0.69 1.065 0.69 1.115 ;
      POLYGON 0.16 1.085 0.16 0.895 0.09 0.895 0.09 0.275 0.175 0.275 0.175 0.105 0.095 0.105 0.095 0.225 0.04 0.225 0.04 0.945 0.11 0.945 0.11 1.085 ;
      POLYGON 0.43 1.08 0.43 0.775 0.225 0.775 0.225 0.375 0.43 0.375 0.43 0.12 0.38 0.12 0.38 0.325 0.175 0.325 0.175 0.825 0.38 0.825 0.38 1.08 ;
      POLYGON 1.51 1.015 1.51 0.875 1.78 0.875 1.78 0.555 1.645 0.555 1.645 0.375 1.375 0.375 1.375 0.165 1.325 0.165 1.325 0.375 1.12 0.375 1.12 0.585 1.17 0.585 1.17 0.425 1.595 0.425 1.595 0.605 1.73 0.605 1.73 0.825 1.46 0.825 1.46 1.015 ;
      POLYGON 0.7 0.945 0.7 0.775 0.785 0.775 0.785 0.835 0.835 0.835 0.835 0.725 0.65 0.725 0.65 0.945 ;
      POLYGON 1.915 0.855 1.915 0.405 2.305 0.405 2.305 0.595 2.54 0.595 2.54 0.525 2.355 0.525 2.355 0.355 2.32 0.355 2.32 0.18 2.27 0.18 2.27 0.355 1.78 0.355 1.78 0.215 1.73 0.215 1.73 0.405 1.865 0.405 1.865 0.855 ;
      POLYGON 2.455 0.835 2.455 0.695 2.66 0.695 2.66 0.585 2.945 0.585 2.945 0.515 2.66 0.515 2.66 0.425 2.455 0.425 2.455 0.165 2.405 0.165 2.405 0.475 2.61 0.475 2.61 0.645 2.405 0.645 2.405 0.785 2.115 0.785 2.115 0.645 2.065 0.645 2.065 0.835 ;
      POLYGON 0.97 0.805 0.97 0.705 1.31 0.705 1.31 0.495 1.26 0.495 1.26 0.655 0.97 0.655 0.97 0.525 0.75 0.525 0.75 0.325 0.835 0.325 0.835 0.15 1 0.15 1 0.1 0.785 0.1 0.785 0.275 0.7 0.275 0.7 0.575 0.92 0.575 0.92 0.805 ;
      POLYGON 1.04 0.475 1.04 0.225 0.905 0.225 0.905 0.275 0.99 0.275 0.99 0.425 0.82 0.425 0.82 0.475 ;
      POLYGON 1.655 0.315 1.655 0.135 2.03 0.135 2.03 0.085 1.585 0.085 1.585 0.315 ;
      RECT 1.845 0.195 2.07 0.275 ;
    LAYER M2 ;
      RECT 0.33 0.925 1.885 0.975 ;
      RECT 0.04 0.225 1.695 0.275 ;
    LAYER VIA1 ;
      RECT 1.705 0.925 1.835 0.975 ;
      RECT 0.93 0.925 1.06 0.975 ;
      RECT 0.38 0.925 0.43 0.975 ;
      RECT 1.595 0.225 1.645 0.275 ;
      RECT 0.95 0.225 1 0.275 ;
      RECT 0.08 0.225 0.13 0.275 ;
  END
END DFFRPQ_X3M_A12TUL_C35

MACRO BUF_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.77 0.875 0.77 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.95 0.16 0.825 0.33 0.825 0.33 0.585 0.65 0.585 0.65 0.515 0.56 0.515 0.56 0.535 0.28 0.535 0.28 0.775 0.09 0.775 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.825 0.11 0.825 0.11 0.95 ;
  END
END BUF_X3M_A12TUL_C35

MACRO AO21B_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011725 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.66 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011725 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.705 0.635 0.705 0.635 0.495 0.58 0.495 0.58 0.705 0.445 0.705 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02135 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.05375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.835 0.37 0.835 0.37 1.165 0.17 1.165 0.17 0.995 0.1 0.995 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.31 1.115 0.31 0.955 0.28 0.955 0.28 0.825 0.075 0.825 0.075 0.355 0.445 0.355 0.445 0.57 0.495 0.57 0.495 0.305 0.16 0.305 0.16 0.12 0.11 0.12 0.11 0.305 0.025 0.305 0.025 0.875 0.23 0.875 0.23 1.115 ;
  END
END AO21B_X0P7M_A12TUL_C35

MACRO AO21B_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00945 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.66 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00945 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.705 0.635 0.705 0.635 0.495 0.58 0.495 0.58 0.705 0.445 0.705 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.085 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.085 ;
    END
    ANTENNADIFFAREA 0.03875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.91 0.37 0.91 0.37 1.165 0.17 1.165 0.17 1.01 0.1 1.01 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.09 0.295 0.825 0.075 0.825 0.075 0.355 0.445 0.355 0.445 0.495 0.495 0.495 0.495 0.305 0.17 0.305 0.17 0.1 0.1 0.1 0.1 0.305 0.025 0.305 0.025 0.875 0.245 0.875 0.245 1.09 ;
  END
END AO21B_X0P5M_A12TUL_C35

MACRO OA21A1OI2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.0745 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.015 0.565 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.515 0.875 0.515 1.015 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OA21A1OI2_X1M_A12TUL_C35

MACRO AO21A1AI2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.015 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.015 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END AO21A1AI2_X0P7M_A12TUL_C35

MACRO AO21A1AI2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.03875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 1.005 0.64 1.005 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END AO21A1AI2_X0P5M_A12TUL_C35

MACRO AO21A1AI2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.07675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.015 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.015 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END AO21A1AI2_X1M_A12TUL_C35

MACRO INV_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X2M_A12TUL_C35

MACRO INV_X5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.161 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.85 0.375 0.85 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
END INV_X5M_A12TUL_C35

MACRO BUF_X3P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X3P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03185 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.905 0.875 0.905 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.85 0.375 0.85 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.27 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.95 0.16 0.825 0.33 0.825 0.33 0.595 0.695 0.595 0.695 0.615 0.785 0.615 0.785 0.545 0.28 0.545 0.28 0.775 0.09 0.775 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.825 0.11 0.825 0.11 0.95 ;
  END
END BUF_X3P5M_A12TUL_C35

MACRO INV_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X1M_A12TUL_C35

MACRO AOI22BB_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22BB_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.77 0.625 0.77 0.445 0.715 0.445 0.715 0.625 0.58 0.625 0.58 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03185 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.585 0.905 0.325 0.685 0.325 0.685 0.375 0.85 0.375 0.85 0.585 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03185 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.615 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B0N
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.705 0.23 0.705 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.915 0.565 0.775 1.04 0.775 1.04 0.225 0.71 0.225 0.71 0.095 0.64 0.095 0.64 0.275 0.985 0.275 0.985 0.725 0.515 0.725 0.515 0.915 ;
    END
    ANTENNADIFFAREA 0.077 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.17 1.165 0.17 0.855 0.1 0.855 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.27 0.575 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.215 0.17 0.215 0.17 0.035 0.37 0.035 0.37 0.215 0.44 0.215 0.44 0.035 0.505 0.035 0.505 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.05 0.43 0.905 0.465 0.905 0.465 0.555 0.65 0.555 0.65 0.485 0.465 0.485 0.465 0.305 0.305 0.305 0.305 0.085 0.235 0.085 0.235 0.355 0.415 0.355 0.415 0.855 0.38 0.855 0.38 1.05 ;
      POLYGON 0.97 1.015 0.97 0.825 0.65 0.825 0.65 1.015 0.7 1.015 0.7 0.875 0.92 0.875 0.92 1.015 ;
  END
END AOI22BB_X1M_A12TUL_C35

MACRO INV_X0P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.07 0.295 0.925 0.365 0.925 0.365 0.09 0.23 0.09 0.23 0.17 0.31 0.17 0.31 0.875 0.245 0.875 0.245 1.07 ;
    END
    ANTENNADIFFAREA 0.028125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.885 0.1 0.885 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.175 0.165 0.175 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.095 0.035 0.095 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P5B_A12TUL_C35

MACRO INV_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X4M_A12TUL_C35

MACRO INV_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X3M_A12TUL_C35

MACRO INV_X3P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X3P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1134 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X3P5M_A12TUL_C35

MACRO BUF_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.025 0.16 0.825 0.33 0.825 0.33 0.595 0.515 0.595 0.515 0.525 0.425 0.525 0.425 0.535 0.28 0.535 0.28 0.775 0.09 0.775 0.09 0.305 0.16 0.305 0.16 0.115 0.11 0.115 0.11 0.255 0.04 0.255 0.04 0.825 0.11 0.825 0.11 1.025 ;
  END
END BUF_X2M_A12TUL_C35

MACRO BUFH_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.595 0.515 0.595 0.515 0.525 0.425 0.525 0.425 0.535 0.28 0.535 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X2M_A12TUL_C35

MACRO BUF_X6M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X6M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05355 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.88 0.785 0.88 0.785 1 0.835 1 0.835 0.88 1.055 0.88 1.055 1 1.105 1 1.105 0.88 1.31 0.88 1.31 0.325 1.105 0.325 1.105 0.205 1.055 0.205 1.055 0.325 0.835 0.325 0.835 0.205 0.785 0.205 0.785 0.325 0.565 0.325 0.565 0.19 0.515 0.19 0.515 0.38 1.255 0.38 1.255 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.27 1.25 0.27 1.25 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 1.1 0.565 1.1 0.585 1.19 0.585 1.19 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUF_X6M_A12TUL_C35

MACRO NAND2_X1B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.07575 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X1B_A12TUL_C35

MACRO XOR3_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.97 0.425 2.02 0.475 ;
        RECT 2.345 0.425 2.395 0.475 ;
      LAYER M1 ;
        RECT 2.335 0.335 2.405 0.625 ;
        POLYGON 1.99 0.635 1.99 0.495 2.07 0.495 2.07 0.425 1.92 0.425 1.92 0.635 ;
      LAYER M2 ;
        RECT 1.92 0.425 2.445 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01995 LAYER M1 ;
    ANTENNAGATEAREA 0.045675 LAYER M2 ;
    ANTENNAGATEAREA 0.045675 LAYER M3 ;
    ANTENNAGATEAREA 0.045675 LAYER M4 ;
    ANTENNAGATEAREA 0.045675 LAYER M5 ;
    ANTENNAGATEAREA 0.045675 LAYER M6 ;
    ANTENNAGATEAREA 0.045675 LAYER M7 ;
    ANTENNAGATEAREA 0.045675 LAYER M8 ;
    ANTENNAGATEAREA 0.045675 LAYER AP ;
    ANTENNAMAXAREACAR 1.017544 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1253133 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.425 0.28 0.425 0.28 0.275 0.715 0.275 0.715 0.135 1.08 0.135 1.08 0.085 0.665 0.085 0.665 0.225 0.23 0.225 0.23 0.375 0.175 0.375 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048125 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.445 0.675 1.445 0.425 1.225 0.425 1.225 0.495 1.39 0.495 1.39 0.625 1.225 0.625 1.225 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04585 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.59 1.015 2.59 0.875 2.795 0.875 2.795 0.325 2.59 0.325 2.59 0.185 2.54 0.185 2.54 0.375 2.74 0.375 2.74 0.825 2.54 0.825 2.54 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
      LAYER M1 ;
        POLYGON 2.835 1.235 2.835 1.165 2.735 1.165 2.735 0.93 2.665 0.93 2.665 1.165 2.47 1.165 2.47 1.03 2.39 1.03 2.39 1.165 1.525 1.165 1.525 1.045 1.445 1.045 1.445 1.165 1.255 1.165 1.255 1.03 1.175 1.03 1.175 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.8 0.235 0.8 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.835 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
      LAYER M1 ;
        POLYGON 2.735 0.27 2.735 0.035 2.835 0.035 2.835 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.525 0.035 0.525 0.12 0.485 0.12 0.485 0.17 0.595 0.17 0.595 0.035 1.16 0.035 1.16 0.165 1.27 0.165 1.27 0.115 1.23 0.115 1.23 0.035 1.445 0.035 1.445 0.155 1.525 0.155 1.525 0.035 2.395 0.035 2.395 0.265 2.465 0.265 2.465 0.035 2.665 0.035 2.665 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 2.835 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.105 1.115 1.105 0.975 1.525 0.975 1.525 0.815 1.575 0.815 1.575 0.325 1.525 0.325 1.525 0.22 0.905 0.22 0.905 0.3 0.985 0.3 0.985 0.27 1.475 0.27 1.475 0.375 1.525 0.375 1.525 0.765 1.475 0.765 1.475 0.925 1.055 0.925 1.055 1.065 0.835 1.065 0.835 0.925 0.785 0.925 0.785 1.115 ;
      POLYGON 1.915 1.065 1.915 0.875 1.71 0.875 1.71 0.27 1.8 0.27 1.8 0.2 1.655 0.2 1.655 0.09 1.585 0.09 1.585 0.27 1.66 0.27 1.66 0.875 1.595 0.875 1.595 1.065 1.645 1.065 1.645 0.925 1.865 0.925 1.865 1.065 ;
      POLYGON 0.16 1.015 0.16 0.725 0.565 0.725 0.565 0.675 0.9 0.675 0.9 0.505 0.85 0.505 0.85 0.625 0.515 0.625 0.515 0.675 0.09 0.675 0.09 0.305 0.16 0.305 0.16 0.115 0.11 0.115 0.11 0.255 0.04 0.255 0.04 0.725 0.11 0.725 0.11 1.015 ;
      POLYGON 0.98 1.005 0.98 0.875 1.405 0.875 1.405 0.825 1.105 0.825 1.105 0.37 1.405 0.37 1.405 0.32 1.055 0.32 1.055 0.825 0.91 0.825 0.91 1.005 ;
      POLYGON 0.43 1 0.43 0.86 0.65 0.86 0.65 0.915 0.7 0.915 0.7 0.775 1.005 0.775 1.005 0.385 0.835 0.385 0.835 0.245 0.785 0.245 0.785 0.325 0.35 0.325 0.35 0.375 0.785 0.375 0.785 0.435 0.955 0.435 0.955 0.725 0.65 0.725 0.65 0.81 0.38 0.81 0.38 1 ;
      POLYGON 2.455 0.975 2.455 0.755 2.52 0.755 2.52 0.575 2.675 0.575 2.675 0.505 2.47 0.505 2.47 0.705 2.405 0.705 2.405 0.925 2.05 0.925 2.05 0.755 1.85 0.755 1.85 0.375 1.925 0.375 1.925 0.195 1.855 0.195 1.855 0.325 1.8 0.325 1.8 0.805 2 0.805 2 0.975 ;
      POLYGON 2.33 0.865 2.33 0.685 2.285 0.685 2.285 0.275 2.32 0.275 2.32 0.085 1.755 0.085 1.755 0.135 2.27 0.135 2.27 0.225 2.235 0.225 2.235 0.73 2.26 0.73 2.26 0.865 ;
      POLYGON 2.185 0.865 2.185 0.325 2.06 0.325 2.06 0.195 1.99 0.195 1.99 0.375 2.135 0.375 2.135 0.865 ;
      RECT 0.29 0.505 0.605 0.575 ;
    LAYER M2 ;
      RECT 1.475 0.725 2.235 0.775 ;
      RECT 0.375 0.525 1.155 0.575 ;
    LAYER VIA1 ;
      RECT 2.135 0.725 2.185 0.775 ;
      RECT 1.525 0.725 1.575 0.775 ;
      RECT 1.055 0.525 1.105 0.575 ;
      RECT 0.425 0.525 0.555 0.575 ;
  END
END XOR3_X2M_A12TUL_C35

MACRO XNOR3_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.85 0.605 1.85 0.295 1.645 0.295 1.645 0.085 1.215 0.085 1.215 0.135 1.595 0.135 1.595 0.345 1.795 0.345 1.795 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.050575 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.805 0.23 0.575 0.58 0.575 0.58 0.715 0.635 0.715 0.635 0.525 0.175 0.525 0.175 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.038325 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.85 0.495 0.85 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.52 1.005 1.52 0.825 1.31 0.825 1.31 0.445 1.375 0.445 1.375 0.255 1.325 0.255 1.325 0.395 1.255 0.395 1.255 0.875 1.45 0.875 1.45 1.005 ;
    END
    ANTENNADIFFAREA 0.08025 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.905 0.235 0.905 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.24 1.79 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.23 0.035 0.23 0.24 0.31 0.24 0.31 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.72 0.035 1.72 0.24 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.645 1.115 1.645 0.875 1.715 0.875 1.715 0.505 1.665 0.505 1.665 0.825 1.595 0.825 1.595 1.065 1.375 1.065 1.375 0.925 1.17 0.925 1.17 0.305 1.255 0.305 1.255 0.225 1.115 0.225 1.115 0.095 1.045 0.095 1.045 0.275 1.12 0.275 1.12 0.925 1.045 0.925 1.045 1.105 1.115 1.105 1.115 0.975 1.325 0.975 1.325 1.115 ;
      POLYGON 0.85 1.115 0.85 0.875 1.04 0.875 1.04 0.325 0.985 0.325 0.985 0.225 0.72 0.225 0.72 0.205 0.63 0.205 0.63 0.275 0.935 0.275 0.935 0.375 0.99 0.375 0.99 0.825 0.8 0.825 0.8 1.065 0.565 1.065 0.565 0.9 0.515 0.9 0.515 1.115 ;
      POLYGON 0.16 1.065 0.16 0.875 0.09 0.875 0.09 0.345 0.43 0.345 0.43 0.135 0.8 0.135 0.8 0.085 0.38 0.085 0.38 0.295 0.16 0.295 0.16 0.235 0.11 0.235 0.11 0.295 0.04 0.295 0.04 0.925 0.11 0.925 0.11 1.065 ;
      POLYGON 0.7 0.995 0.7 0.835 0.74 0.835 0.74 0.775 0.865 0.775 0.865 0.725 0.74 0.725 0.74 0.375 0.865 0.375 0.865 0.325 0.69 0.325 0.69 0.785 0.365 0.785 0.365 0.635 0.315 0.635 0.315 0.835 0.65 0.835 0.65 0.995 ;
      POLYGON 1.915 0.945 1.915 0.785 1.98 0.785 1.98 0.175 1.845 0.175 1.845 0.245 1.93 0.245 1.93 0.715 1.775 0.715 1.775 0.785 1.865 0.785 1.865 0.945 ;
      POLYGON 1.605 0.775 1.605 0.705 1.44 0.705 1.44 0.515 1.39 0.515 1.39 0.775 ;
      POLYGON 0.565 0.455 0.565 0.265 0.515 0.265 0.515 0.405 0.35 0.405 0.35 0.455 ;
      POLYGON 1.675 0.445 1.675 0.395 1.51 0.395 1.51 0.255 1.46 0.255 1.46 0.445 ;
    LAYER M2 ;
      RECT 1.465 0.725 1.985 0.775 ;
    LAYER VIA1 ;
      RECT 1.805 0.725 1.935 0.775 ;
      RECT 1.515 0.725 1.565 0.775 ;
  END
END XNOR3_X1M_A12TUL_C35

MACRO BUF_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0364 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.85 0.1 0.85 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.025 0.295 0.775 0.495 0.775 0.495 0.565 0.83 0.565 0.83 0.585 0.92 0.585 0.92 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.115 0.245 0.115 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 1.025 ;
  END
END BUF_X4M_A12TUL_C35

MACRO XOR3_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.85 0.605 1.85 0.295 1.645 0.295 1.645 0.085 1.21 0.085 1.21 0.135 1.595 0.135 1.595 0.345 1.795 0.345 1.795 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.050575 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.805 0.23 0.575 0.58 0.575 0.58 0.715 0.635 0.715 0.635 0.525 0.175 0.525 0.175 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03885 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.705 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.845 0.495 0.845 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.52 1.005 1.52 0.825 1.31 0.825 1.31 0.445 1.375 0.445 1.375 0.255 1.325 0.255 1.325 0.395 1.255 0.395 1.255 0.875 1.45 0.875 1.45 1.005 ;
    END
    ANTENNADIFFAREA 0.080625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 0.985 1.165 0.985 1.055 0.905 1.055 0.905 1.165 0.305 1.165 0.305 0.905 0.235 0.905 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.375 0.305 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.72 0.035 1.72 0.24 1.79 0.24 1.79 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.645 1.115 1.645 0.875 1.715 0.875 1.715 0.505 1.665 0.505 1.665 0.825 1.595 0.825 1.595 1.065 1.375 1.065 1.375 0.925 1.17 0.925 1.17 0.3 1.255 0.3 1.255 0.22 1.115 0.22 1.115 0.09 1.045 0.09 1.045 0.27 1.12 0.27 1.12 0.925 1.045 0.925 1.045 1.105 1.115 1.105 1.115 0.975 1.325 0.975 1.325 1.115 ;
      POLYGON 0.835 1.095 0.835 1.005 0.97 1.005 0.97 0.84 1.035 0.84 1.035 0.325 0.985 0.325 0.985 0.225 0.515 0.225 0.515 0.415 0.565 0.415 0.565 0.275 0.935 0.275 0.935 0.375 0.985 0.375 0.985 0.79 0.92 0.79 0.92 0.955 0.785 0.955 0.785 1.045 0.7 1.045 0.7 0.905 0.65 0.905 0.65 1.095 ;
      POLYGON 0.565 1.085 0.565 0.895 0.38 0.895 0.38 1.085 0.43 1.085 0.43 0.945 0.515 0.945 0.515 1.085 ;
      POLYGON 0.16 1.065 0.16 0.875 0.09 0.875 0.09 0.475 0.43 0.475 0.43 0.135 0.795 0.135 0.795 0.085 0.38 0.085 0.38 0.425 0.16 0.425 0.16 0.365 0.11 0.365 0.11 0.425 0.04 0.425 0.04 0.925 0.11 0.925 0.11 1.065 ;
      POLYGON 1.915 0.945 1.915 0.785 1.98 0.785 1.98 0.175 1.845 0.175 1.845 0.245 1.93 0.245 1.93 0.715 1.775 0.715 1.775 0.785 1.865 0.785 1.865 0.945 ;
      POLYGON 0.85 0.905 0.85 0.785 0.76 0.785 0.76 0.375 0.865 0.375 0.865 0.325 0.635 0.325 0.635 0.4 0.71 0.4 0.71 0.785 0.36 0.785 0.36 0.675 0.31 0.675 0.31 0.835 0.77 0.835 0.77 0.905 ;
      POLYGON 1.605 0.775 1.605 0.705 1.44 0.705 1.44 0.515 1.39 0.515 1.39 0.775 ;
      POLYGON 1.675 0.445 1.675 0.395 1.51 0.395 1.51 0.255 1.46 0.255 1.46 0.445 ;
    LAYER M2 ;
      RECT 1.465 0.725 1.985 0.775 ;
    LAYER VIA1 ;
      RECT 1.805 0.725 1.935 0.775 ;
      RECT 1.515 0.725 1.565 0.775 ;
  END
END XOR3_X1M_A12TUL_C35

MACRO XOR3_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.295 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.28 0.925 0.33 0.975 ;
        RECT 1.215 0.925 1.345 0.975 ;
      LAYER M1 ;
        POLYGON 0.36 0.975 0.36 0.63 0.31 0.63 0.31 0.905 0.25 0.905 0.25 0.975 ;
        POLYGON 1.605 1.075 1.605 1.025 1.385 1.025 1.385 0.925 1.175 0.925 1.175 0.975 1.335 0.975 1.335 1.075 ;
      LAYER M2 ;
        RECT 0.23 0.925 1.395 0.975 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 LAYER M1 ;
    ANTENNAGATEAREA 0.04025 LAYER M2 ;
    ANTENNAGATEAREA 0.04025 LAYER M3 ;
    ANTENNAGATEAREA 0.04025 LAYER M4 ;
    ANTENNAGATEAREA 0.04025 LAYER M5 ;
    ANTENNAGATEAREA 0.04025 LAYER M6 ;
    ANTENNAGATEAREA 0.04025 LAYER M7 ;
    ANTENNAGATEAREA 0.04025 LAYER M8 ;
    ANTENNAGATEAREA 0.04025 LAYER AP ;
    ANTENNAMAXAREACAR 1.459184 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4421769 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.19 0.525 0.24 0.575 ;
        RECT 1.135 0.525 1.185 0.575 ;
      LAYER M1 ;
        RECT 1.12 0.455 1.205 0.645 ;
        RECT 0.18 0.41 0.25 0.725 ;
      LAYER M2 ;
        RECT 0.14 0.525 1.235 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 LAYER M1 ;
    ANTENNAGATEAREA 0.05075 LAYER M2 ;
    ANTENNAGATEAREA 0.05075 LAYER M3 ;
    ANTENNAGATEAREA 0.05075 LAYER M4 ;
    ANTENNAGATEAREA 0.05075 LAYER M5 ;
    ANTENNAGATEAREA 0.05075 LAYER M6 ;
    ANTENNAGATEAREA 0.05075 LAYER M7 ;
    ANTENNAGATEAREA 0.05075 LAYER M8 ;
    ANTENNAGATEAREA 0.05075 LAYER AP ;
    ANTENNAMAXAREACAR 1.166667 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1322753 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.565 0.295 0.635 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03115 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.05 1.105 2.05 0.965 2.085 0.965 2.085 0.875 2.255 0.875 2.255 0.325 2.05 0.325 2.05 0.175 2 0.175 2 0.375 2.2 0.375 2.2 0.825 2.035 0.825 2.035 0.915 2 0.915 2 1.105 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
      LAYER M1 ;
        POLYGON 2.295 1.235 2.295 1.165 2.205 1.165 2.205 0.925 2.135 0.925 2.135 1.165 1.93 1.165 1.93 0.955 1.85 0.955 1.85 1.165 0.715 1.165 0.715 0.96 0.635 0.96 0.635 1.165 0.305 1.165 0.305 1.04 0.235 1.04 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.295 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.31 0.305 0.035 0.635 0.035 0.635 0.145 0.715 0.145 0.715 0.035 1.855 0.035 1.855 0.16 1.925 0.16 1.925 0.035 2.125 0.035 2.125 0.27 2.195 0.27 2.195 0.035 2.295 0.035 2.295 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.31 ;
      LAYER M2 ;
        RECT 0 -0.065 2.295 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.46 1.105 0.46 0.475 0.43 0.475 0.43 0.095 0.38 0.095 0.38 0.525 0.41 0.525 0.41 1.025 0.365 1.025 0.365 1.105 ;
      POLYGON 0.97 1.045 0.97 0.855 0.735 0.855 0.735 0.595 0.785 0.595 0.785 0.525 0.735 0.525 0.735 0.245 0.85 0.245 0.85 0.135 1.19 0.135 1.19 0.275 1.24 0.275 1.24 0.085 0.8 0.085 0.8 0.195 0.58 0.195 0.58 0.165 0.5 0.165 0.5 0.245 0.685 0.245 0.685 0.855 0.515 0.855 0.515 1.045 0.565 1.045 0.565 0.905 0.92 0.905 0.92 1.045 ;
      POLYGON 0.16 1.035 0.16 0.845 0.13 0.845 0.13 0.325 0.16 0.325 0.16 0.135 0.11 0.135 0.11 0.275 0.08 0.275 0.08 0.895 0.11 0.895 0.11 1.035 ;
      POLYGON 1.105 1.015 1.105 0.875 1.375 0.875 1.375 0.595 1.34 0.595 1.34 0.275 1.52 0.275 1.52 0.095 1.45 0.095 1.45 0.225 1.29 0.225 1.29 0.345 1.105 0.345 1.105 0.205 1.055 0.205 1.055 0.395 1.29 0.395 1.29 0.645 1.325 0.645 1.325 0.825 1.055 0.825 1.055 1.015 ;
      POLYGON 1.915 0.905 1.915 0.855 1.985 0.855 1.985 0.475 2.065 0.475 2.065 0.615 2.115 0.615 2.115 0.425 1.94 0.425 1.94 0.225 1.655 0.225 1.655 0.095 1.585 0.095 1.585 0.275 1.89 0.275 1.89 0.475 1.935 0.475 1.935 0.805 1.865 0.805 1.865 0.855 1.525 0.855 1.525 0.745 1.445 0.745 1.445 0.905 ;
      POLYGON 1.78 0.8 1.78 0.69 1.73 0.69 1.73 0.75 1.66 0.75 1.66 0.64 1.58 0.64 1.58 0.375 1.82 0.375 1.82 0.325 1.53 0.325 1.53 0.69 1.58 0.69 1.58 0.8 ;
      RECT 0.785 0.665 0.89 0.775 ;
      POLYGON 1.26 0.775 1.26 0.705 1.17 0.705 1.17 0.725 0.89 0.725 0.89 0.455 0.97 0.455 0.97 0.265 0.92 0.265 0.92 0.405 0.835 0.405 0.835 0.315 0.785 0.315 0.785 0.455 0.84 0.455 0.84 0.665 0.785 0.665 0.785 0.775 ;
      POLYGON 1.885 0.735 1.885 0.525 1.78 0.525 1.78 0.605 1.83 0.605 1.83 0.735 ;
      POLYGON 1.055 0.675 1.055 0.505 0.975 0.505 0.975 0.605 0.945 0.605 0.945 0.675 ;
      POLYGON 1.72 0.585 1.72 0.475 1.79 0.475 1.79 0.425 1.64 0.425 1.64 0.585 ;
      RECT 1.39 0.33 1.465 0.54 ;
    LAYER M2 ;
      RECT 1.275 0.625 1.935 0.675 ;
      RECT 0.04 0.625 1.075 0.675 ;
      RECT 0.33 0.425 1.79 0.475 ;
    LAYER VIA1 ;
      RECT 1.835 0.625 1.885 0.675 ;
      RECT 1.325 0.625 1.375 0.675 ;
      RECT 0.975 0.625 1.025 0.675 ;
      RECT 0.08 0.625 0.13 0.675 ;
      RECT 1.69 0.425 1.74 0.475 ;
      RECT 1.405 0.425 1.455 0.475 ;
      RECT 0.38 0.425 0.43 0.475 ;
  END
END XOR3_X1P4M_A12TUL_C35

MACRO BUF_X5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.215 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0448 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.175 0.875 1.175 0.325 1.105 0.325 1.105 0.2 1.055 0.2 1.055 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 1.12 0.375 1.12 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
      LAYER M1 ;
        POLYGON 1.215 1.235 1.215 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.215 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.215 0.035 1.215 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.215 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.96 0.295 0.775 0.495 0.775 0.495 0.565 0.965 0.565 0.965 0.585 1.055 0.585 1.055 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.17 0.245 0.17 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.96 ;
  END
END BUF_X5M_A12TUL_C35

MACRO INV_X9M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X9M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.575 1.255 0.575 1.255 0.605 1.31 0.605 1.31 0.495 1.255 0.495 1.255 0.525 0.905 0.525 0.905 0.425 0.685 0.425 0.685 0.475 0.855 0.475 0.855 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 0.635 0.675 0.635 0.575 1.125 0.575 1.125 0.625 0.955 0.625 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2898 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.89 0.515 0.89 0.515 0.985 0.565 0.985 0.565 0.89 0.785 0.89 0.785 0.985 0.835 0.985 0.835 0.89 1.055 0.89 1.055 0.985 1.105 0.985 1.105 0.89 1.325 0.89 1.325 0.985 1.375 0.985 1.375 0.89 1.46 0.89 1.46 0.295 1.375 0.295 1.375 0.195 1.325 0.195 1.325 0.295 1.105 0.295 1.105 0.2 1.055 0.2 1.055 0.295 0.835 0.295 0.835 0.2 0.785 0.2 0.785 0.295 0.565 0.295 0.565 0.2 0.515 0.2 0.515 0.295 0.295 0.295 0.295 0.185 0.245 0.185 0.245 0.375 1.38 0.375 1.38 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.437 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 1.255 1.165 1.255 0.955 1.175 0.955 1.175 1.165 0.985 1.165 0.985 0.955 0.905 0.955 0.905 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.365 0.035 0.365 0.235 0.445 0.235 0.445 0.035 0.635 0.035 0.635 0.235 0.715 0.235 0.715 0.035 0.905 0.035 0.905 0.235 0.985 0.235 0.985 0.035 1.175 0.035 1.175 0.235 1.255 0.235 1.255 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
END INV_X9M_A12TUL_C35

MACRO INV_X7P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X7P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.675 1.04 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.77 0.525 0.77 0.425 0.55 0.425 0.55 0.475 0.72 0.475 0.72 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2422 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.88 0.515 0.88 0.515 0.985 0.565 0.985 0.565 0.88 0.785 0.88 0.785 0.985 0.835 0.985 0.835 0.88 1.055 0.88 1.055 0.985 1.105 0.985 1.105 0.88 1.325 0.88 1.325 0.305 1.105 0.305 1.105 0.2 1.055 0.2 1.055 0.305 0.835 0.305 0.835 0.2 0.785 0.2 0.785 0.305 0.565 0.305 0.565 0.2 0.515 0.2 0.515 0.305 0.295 0.305 0.295 0.185 0.245 0.185 0.245 0.375 1.255 0.375 1.255 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.245 0.44 0.245 0.44 0.035 0.64 0.035 0.64 0.245 0.71 0.245 0.71 0.035 0.91 0.035 0.91 0.245 0.98 0.245 0.98 0.035 1.175 0.035 1.175 0.255 1.255 0.255 1.255 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
END INV_X7P5M_A12TUL_C35

MACRO XNOR3_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.645 1.105 1.645 0.675 1.85 0.675 1.85 0.395 1.795 0.395 1.795 0.625 1.58 0.625 1.58 0.495 1.525 0.495 1.525 0.675 1.595 0.675 1.595 1.055 1.23 1.055 1.23 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.041475 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.415 0.475 0.415 0.135 0.795 0.135 0.795 0.085 0.365 0.085 0.365 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03675 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.85 0.495 0.85 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01925 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.525 0.995 1.525 0.825 1.31 0.825 1.31 0.375 1.405 0.375 1.405 0.325 1.255 0.325 1.255 0.875 1.45 0.875 1.45 0.995 ;
    END
    ANTENNADIFFAREA 0.068875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.845 1.72 0.845 1.72 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.72 0.035 1.72 0.29 1.79 0.29 1.79 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.115 1.105 1.115 0.975 1.305 0.975 1.305 0.995 1.395 0.995 1.395 0.925 1.17 0.925 1.17 0.275 1.48 0.275 1.48 0.425 1.66 0.425 1.66 0.505 1.71 0.505 1.71 0.375 1.53 0.375 1.53 0.225 1.24 0.225 1.24 0.1 1.19 0.1 1.19 0.225 1.115 0.225 1.115 0.095 1.045 0.095 1.045 0.275 1.12 0.275 1.12 0.925 1.045 0.925 1.045 1.105 ;
      POLYGON 0.565 1.085 0.565 0.825 0.515 0.825 0.515 1.035 0.43 1.035 0.43 0.895 0.38 0.895 0.38 1.085 ;
      POLYGON 0.16 1.075 0.16 0.825 0.465 0.825 0.465 0.755 0.635 0.755 0.635 0.505 0.585 0.505 0.585 0.705 0.415 0.705 0.415 0.775 0.105 0.775 0.105 0.345 0.175 0.345 0.175 0.265 0.055 0.265 0.055 0.825 0.11 0.825 0.11 1.075 ;
      POLYGON 0.7 1.015 0.7 0.875 1.04 0.875 1.04 0.325 0.985 0.325 0.985 0.225 0.485 0.225 0.485 0.275 0.935 0.275 0.935 0.375 0.99 0.375 0.99 0.825 0.65 0.825 0.65 1.015 ;
      POLYGON 1.915 0.935 1.915 0.775 1.995 0.775 1.995 0.175 1.85 0.175 1.85 0.255 1.945 0.255 1.945 0.725 1.755 0.725 1.755 0.775 1.865 0.775 1.865 0.935 ;
      POLYGON 1.525 0.775 1.525 0.725 1.45 0.725 1.45 0.475 1.38 0.475 1.38 0.775 ;
      POLYGON 0.865 0.775 0.865 0.725 0.75 0.725 0.75 0.375 0.865 0.375 0.865 0.325 0.475 0.325 0.475 0.525 0.3 0.525 0.3 0.7 0.36 0.7 0.36 0.575 0.525 0.575 0.525 0.375 0.7 0.375 0.7 0.775 ;
      POLYGON 1.645 0.3 1.645 0.11 1.43 0.11 1.43 0.16 1.595 0.16 1.595 0.3 ;
    LAYER M2 ;
      RECT 1.375 0.725 1.985 0.775 ;
    LAYER VIA1 ;
      RECT 1.805 0.725 1.935 0.775 ;
      RECT 1.425 0.725 1.475 0.775 ;
  END
END XNOR3_X0P7M_A12TUL_C35

MACRO XNOR3_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.85 0.605 1.85 0.345 1.795 0.345 1.795 0.295 1.645 0.295 1.645 0.085 1.23 0.085 1.23 0.135 1.595 0.135 1.595 0.345 1.745 0.345 1.745 0.395 1.795 0.395 1.795 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.415 0.475 0.415 0.155 0.795 0.155 0.795 0.105 0.365 0.105 0.365 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.028 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.85 0.495 0.85 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0161 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.525 1.01 1.525 0.825 1.31 0.825 1.31 0.445 1.375 0.445 1.375 0.255 1.325 0.255 1.325 0.395 1.255 0.395 1.255 0.875 1.445 0.875 1.445 1.01 ;
    END
    ANTENNADIFFAREA 0.05875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.885 1.72 0.885 1.72 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.905 0.235 0.905 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.31 0.375 0.31 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.715 0.035 1.715 0.245 1.795 0.245 1.795 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.23 0.035 0.23 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.645 1.115 1.645 0.815 1.74 0.815 1.74 0.765 1.595 0.765 1.595 1.065 1.375 1.065 1.375 0.925 1.17 0.925 1.17 0.3 1.255 0.3 1.255 0.22 1.115 0.22 1.115 0.09 1.045 0.09 1.045 0.27 1.12 0.27 1.12 0.925 1.045 0.925 1.045 1.105 1.115 1.105 1.115 0.975 1.325 0.975 1.325 1.115 ;
      POLYGON 0.43 1.095 0.43 0.955 0.565 0.955 0.565 0.755 0.515 0.755 0.515 0.905 0.38 0.905 0.38 1.095 ;
      POLYGON 0.16 1.07 0.16 0.835 0.465 0.835 0.465 0.685 0.635 0.685 0.635 0.505 0.585 0.505 0.585 0.635 0.415 0.635 0.415 0.785 0.09 0.785 0.09 0.315 0.175 0.315 0.175 0.235 0.04 0.235 0.04 0.835 0.11 0.835 0.11 1.07 ;
      POLYGON 1.915 1.035 1.915 0.715 1.985 0.715 1.985 0.2 1.85 0.2 1.85 0.28 1.935 0.28 1.935 0.665 1.44 0.665 1.44 0.525 1.39 0.525 1.39 0.715 1.865 0.715 1.865 1.035 ;
      POLYGON 0.72 0.895 0.72 0.875 1.035 0.875 1.035 0.325 0.985 0.325 0.985 0.225 0.485 0.225 0.485 0.275 0.935 0.275 0.935 0.375 0.985 0.375 0.985 0.825 0.63 0.825 0.63 0.895 ;
      POLYGON 0.865 0.775 0.865 0.725 0.75 0.725 0.75 0.375 0.865 0.375 0.865 0.325 0.475 0.325 0.475 0.525 0.31 0.525 0.31 0.715 0.36 0.715 0.36 0.575 0.525 0.575 0.525 0.375 0.7 0.375 0.7 0.775 ;
      POLYGON 1.675 0.445 1.675 0.395 1.51 0.395 1.51 0.255 1.46 0.255 1.46 0.445 ;
  END
END XNOR3_X0P5M_A12TUL_C35

MACRO INV_X6M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X6M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.5 0.525 0.5 0.425 0.28 0.425 0.28 0.475 0.45 0.475 0.45 0.525 0.145 0.525 0.145 0.575 0.72 0.575 0.72 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1932 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.01 0.295 0.875 0.515 0.875 0.515 0.995 0.565 0.995 0.565 0.875 0.785 0.875 0.785 0.995 0.835 0.995 0.835 0.875 1.04 0.875 1.04 0.32 0.835 0.32 0.835 0.2 0.785 0.2 0.785 0.32 0.565 0.32 0.565 0.2 0.515 0.2 0.515 0.32 0.295 0.32 0.295 0.185 0.245 0.185 0.245 0.375 0.985 0.375 0.985 0.82 0.245 0.82 0.245 1.01 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
END INV_X6M_A12TUL_C35

MACRO BUF_X7P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X7P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.995 0.565 0.875 0.785 0.875 0.785 0.98 0.835 0.98 0.835 0.875 1.055 0.875 1.055 0.98 1.105 0.98 1.105 0.875 1.325 0.875 1.325 0.98 1.375 0.98 1.375 0.875 1.585 0.875 1.585 0.325 1.375 0.325 1.375 0.22 1.325 0.22 1.325 0.325 1.105 0.325 1.105 0.22 1.055 0.22 1.055 0.325 0.835 0.325 0.835 0.22 0.785 0.22 0.785 0.325 0.565 0.325 0.565 0.205 0.515 0.205 0.515 0.395 1.515 0.395 1.515 0.805 0.515 0.805 0.515 0.995 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 1.52 1.165 1.52 0.93 1.45 0.93 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.27 1.52 0.27 1.52 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.43 0.775 0.43 0.725 0.5 0.725 0.5 0.56 1.375 0.56 1.375 0.6 1.455 0.6 1.455 0.51 0.45 0.51 0.45 0.675 0.38 0.675 0.38 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUF_X7P5M_A12TUL_C35

MACRO XNOR3_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.295 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.28 0.925 0.33 0.975 ;
        RECT 1.215 0.925 1.345 0.975 ;
      LAYER M1 ;
        POLYGON 0.36 0.975 0.36 0.63 0.31 0.63 0.31 0.905 0.25 0.905 0.25 0.975 ;
        POLYGON 1.605 1.075 1.605 1.025 1.385 1.025 1.385 0.925 1.175 0.925 1.175 0.975 1.335 0.975 1.335 1.075 ;
      LAYER M2 ;
        RECT 0.23 0.925 1.395 0.975 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 LAYER M1 ;
    ANTENNAGATEAREA 0.04025 LAYER M2 ;
    ANTENNAGATEAREA 0.04025 LAYER M3 ;
    ANTENNAGATEAREA 0.04025 LAYER M4 ;
    ANTENNAGATEAREA 0.04025 LAYER M5 ;
    ANTENNAGATEAREA 0.04025 LAYER M6 ;
    ANTENNAGATEAREA 0.04025 LAYER M7 ;
    ANTENNAGATEAREA 0.04025 LAYER M8 ;
    ANTENNAGATEAREA 0.04025 LAYER AP ;
    ANTENNAMAXAREACAR 1.459184 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4421769 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.19 0.625 0.24 0.675 ;
        RECT 0.975 0.625 1.025 0.675 ;
      LAYER M1 ;
        POLYGON 1.055 0.675 1.055 0.505 0.975 0.505 0.975 0.605 0.945 0.605 0.945 0.675 ;
        RECT 0.18 0.41 0.25 0.725 ;
      LAYER M2 ;
        RECT 0.14 0.625 1.075 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 LAYER M1 ;
    ANTENNAGATEAREA 0.05075 LAYER M2 ;
    ANTENNAGATEAREA 0.05075 LAYER M3 ;
    ANTENNAGATEAREA 0.05075 LAYER M4 ;
    ANTENNAGATEAREA 0.05075 LAYER M5 ;
    ANTENNAGATEAREA 0.05075 LAYER M6 ;
    ANTENNAGATEAREA 0.05075 LAYER M7 ;
    ANTENNAGATEAREA 0.05075 LAYER M8 ;
    ANTENNAGATEAREA 0.05075 LAYER AP ;
    ANTENNAMAXAREACAR 1.166667 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1322753 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.565 0.295 0.635 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03115 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.05 1.105 2.05 0.965 2.085 0.965 2.085 0.875 2.255 0.875 2.255 0.325 2.05 0.325 2.05 0.175 2 0.175 2 0.375 2.2 0.375 2.2 0.825 2.035 0.825 2.035 0.915 2 0.915 2 1.105 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
      LAYER M1 ;
        POLYGON 2.295 1.235 2.295 1.165 2.205 1.165 2.205 0.925 2.135 0.925 2.135 1.165 1.93 1.165 1.93 0.955 1.85 0.955 1.85 1.165 0.715 1.165 0.715 0.96 0.635 0.96 0.635 1.165 0.305 1.165 0.305 1.04 0.235 1.04 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.295 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.31 0.305 0.035 0.635 0.035 0.635 0.145 0.715 0.145 0.715 0.035 1.855 0.035 1.855 0.16 1.925 0.16 1.925 0.035 2.125 0.035 2.125 0.27 2.195 0.27 2.195 0.035 2.295 0.035 2.295 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.31 ;
      LAYER M2 ;
        RECT 0 -0.065 2.295 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.46 1.105 0.46 0.475 0.43 0.475 0.43 0.095 0.38 0.095 0.38 0.525 0.41 0.525 0.41 1.025 0.365 1.025 0.365 1.105 ;
      POLYGON 0.97 1.045 0.97 0.855 0.735 0.855 0.735 0.595 0.785 0.595 0.785 0.525 0.735 0.525 0.735 0.245 0.85 0.245 0.85 0.135 1.19 0.135 1.19 0.275 1.24 0.275 1.24 0.085 0.8 0.085 0.8 0.195 0.58 0.195 0.58 0.165 0.5 0.165 0.5 0.245 0.685 0.245 0.685 0.855 0.515 0.855 0.515 1.045 0.565 1.045 0.565 0.905 0.92 0.905 0.92 1.045 ;
      POLYGON 0.16 1.035 0.16 0.845 0.13 0.845 0.13 0.325 0.16 0.325 0.16 0.135 0.11 0.135 0.11 0.275 0.08 0.275 0.08 0.895 0.11 0.895 0.11 1.035 ;
      POLYGON 1.105 1.015 1.105 0.875 1.375 0.875 1.375 0.595 1.34 0.595 1.34 0.275 1.52 0.275 1.52 0.095 1.45 0.095 1.45 0.225 1.29 0.225 1.29 0.345 1.105 0.345 1.105 0.205 1.055 0.205 1.055 0.395 1.29 0.395 1.29 0.645 1.325 0.645 1.325 0.825 1.055 0.825 1.055 1.015 ;
      POLYGON 1.915 0.905 1.915 0.855 1.985 0.855 1.985 0.475 2.065 0.475 2.065 0.615 2.115 0.615 2.115 0.425 1.94 0.425 1.94 0.225 1.655 0.225 1.655 0.095 1.585 0.095 1.585 0.275 1.89 0.275 1.89 0.475 1.935 0.475 1.935 0.805 1.865 0.805 1.865 0.855 1.525 0.855 1.525 0.745 1.445 0.745 1.445 0.905 ;
      POLYGON 1.78 0.8 1.78 0.69 1.73 0.69 1.73 0.75 1.66 0.75 1.66 0.64 1.58 0.64 1.58 0.375 1.82 0.375 1.82 0.325 1.53 0.325 1.53 0.69 1.58 0.69 1.58 0.8 ;
      RECT 0.785 0.665 0.89 0.775 ;
      POLYGON 1.26 0.775 1.26 0.705 1.17 0.705 1.17 0.725 0.89 0.725 0.89 0.455 0.97 0.455 0.97 0.265 0.92 0.265 0.92 0.405 0.835 0.405 0.835 0.315 0.785 0.315 0.785 0.455 0.84 0.455 0.84 0.665 0.785 0.665 0.785 0.775 ;
      POLYGON 1.885 0.735 1.885 0.525 1.78 0.525 1.78 0.605 1.83 0.605 1.83 0.735 ;
      RECT 1.12 0.455 1.205 0.645 ;
      POLYGON 1.72 0.585 1.72 0.475 1.79 0.475 1.79 0.425 1.64 0.425 1.64 0.585 ;
      RECT 1.39 0.33 1.465 0.54 ;
    LAYER M2 ;
      RECT 1.275 0.625 1.935 0.675 ;
      RECT 0.04 0.525 1.235 0.575 ;
      RECT 0.33 0.425 1.79 0.475 ;
    LAYER VIA1 ;
      RECT 1.835 0.625 1.885 0.675 ;
      RECT 1.325 0.625 1.375 0.675 ;
      RECT 1.135 0.525 1.185 0.575 ;
      RECT 0.08 0.525 0.13 0.575 ;
      RECT 1.69 0.425 1.74 0.475 ;
      RECT 1.405 0.425 1.455 0.475 ;
      RECT 0.38 0.425 0.43 0.475 ;
  END
END XNOR3_X1P4M_A12TUL_C35

MACRO BUFH_X11M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X11M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.635 0.525 0.635 0.425 0.415 0.425 0.415 0.475 0.585 0.475 0.585 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 0.365 0.675 0.365 0.575 0.72 0.575 0.72 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1932 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.105 0.98 1.105 0.885 1.325 0.885 1.325 0.965 1.375 0.965 1.375 0.885 1.595 0.885 1.595 0.965 1.645 0.965 1.645 0.885 1.865 0.885 1.865 0.965 1.915 0.965 1.915 0.885 2.135 0.885 2.135 0.965 2.185 0.965 2.185 0.885 2.405 0.885 2.405 0.965 2.455 0.965 2.455 0.885 2.54 0.885 2.54 0.315 2.455 0.315 2.455 0.235 2.405 0.235 2.405 0.315 2.185 0.315 2.185 0.235 2.135 0.235 2.135 0.315 1.915 0.315 1.915 0.235 1.865 0.235 1.865 0.315 1.645 0.315 1.645 0.235 1.595 0.235 1.595 0.315 1.375 0.315 1.375 0.235 1.325 0.235 1.325 0.315 1.105 0.315 1.105 0.22 1.055 0.22 1.055 0.41 2.445 0.41 2.445 0.79 1.055 0.79 1.055 0.98 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
      LAYER M1 ;
        POLYGON 2.565 1.235 2.565 1.165 2.33 1.165 2.33 0.945 2.26 0.945 2.26 1.165 2.06 1.165 2.06 0.945 1.99 0.945 1.99 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.845 0.91 0.845 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.565 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.355 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 1.72 0.035 1.72 0.255 1.79 0.255 1.79 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.26 0.035 2.26 0.255 2.33 0.255 2.33 0.035 2.565 0.035 2.565 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.565 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.835 0.9 0.835 0.775 0.97 0.775 0.97 0.715 1.035 0.715 1.035 0.565 2.325 0.565 2.325 0.605 2.395 0.605 2.395 0.515 0.985 0.515 0.985 0.665 0.92 0.665 0.92 0.725 0.075 0.725 0.075 0.375 0.835 0.375 0.835 0.185 0.785 0.185 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 0.295 0.9 0.295 0.775 0.515 0.775 0.515 0.9 0.565 0.9 0.565 0.775 0.785 0.775 0.785 0.9 ;
  END
END BUFH_X11M_A12TUL_C35

MACRO BUFH_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.525 0.145 0.525 0.145 0.575 0.345 0.575 0.345 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 0.84 0.565 0.84 0.605 0.91 0.605 0.91 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUFH_X4M_A12TUL_C35

MACRO XOR3_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.51 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.795 0.625 1.845 0.675 ;
        RECT 2.785 0.625 2.835 0.675 ;
      LAYER M1 ;
        POLYGON 2.91 0.675 2.91 0.605 2.815 0.605 2.815 0.515 2.735 0.515 2.735 0.675 ;
        RECT 1.785 0.42 1.855 0.71 ;
      LAYER M2 ;
        RECT 1.745 0.625 2.885 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 LAYER M1 ;
    ANTENNAGATEAREA 0.05495 LAYER M2 ;
    ANTENNAGATEAREA 0.05495 LAYER M3 ;
    ANTENNAGATEAREA 0.05495 LAYER M4 ;
    ANTENNAGATEAREA 0.05495 LAYER M5 ;
    ANTENNAGATEAREA 0.05495 LAYER M6 ;
    ANTENNAGATEAREA 0.05495 LAYER M7 ;
    ANTENNAGATEAREA 0.05495 LAYER M8 ;
    ANTENNAGATEAREA 0.05495 LAYER AP ;
    ANTENNAMAXAREACAR 0.8923078 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1098901 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.15 0.525 1.28 0.575 ;
        RECT 1.66 0.525 1.71 0.575 ;
      LAYER M1 ;
        POLYGON 1.32 0.63 1.32 0.515 1.11 0.515 1.11 0.63 1.18 0.63 1.18 0.585 1.25 0.585 1.25 0.63 ;
        RECT 1.65 0.42 1.72 0.71 ;
      LAYER M2 ;
        RECT 1.1 0.525 1.76 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0308 LAYER M1 ;
    ANTENNAGATEAREA 0.0924 LAYER M2 ;
    ANTENNAGATEAREA 0.0924 LAYER M3 ;
    ANTENNAGATEAREA 0.0924 LAYER M4 ;
    ANTENNAGATEAREA 0.0924 LAYER M5 ;
    ANTENNAGATEAREA 0.0924 LAYER M6 ;
    ANTENNAGATEAREA 0.0924 LAYER M7 ;
    ANTENNAGATEAREA 0.0924 LAYER M8 ;
    ANTENNAGATEAREA 0.0924 LAYER AP ;
    ANTENNAMAXAREACAR 0.659091 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.211039 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.465 0.625 0.465 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05775 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 3.13 1.015 3.13 0.875 3.35 0.875 3.35 1 3.4 1 3.4 0.875 3.47 0.875 3.47 0.325 3.4 0.325 3.4 0.19 3.35 0.19 3.35 0.325 3.13 0.325 3.13 0.185 3.08 0.185 3.08 0.375 3.415 0.375 3.415 0.825 3.08 0.825 3.08 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
      LAYER M1 ;
        POLYGON 3.51 1.235 3.51 1.165 3.275 1.165 3.275 0.945 3.205 0.945 3.205 1.165 3.005 1.165 3.005 0.845 2.935 0.845 2.935 1.165 2.47 1.165 2.47 1.03 2.39 1.03 2.39 1.165 2.195 1.165 2.195 0.915 2.125 0.915 2.125 1.165 1.79 1.165 1.79 0.78 1.72 0.78 1.72 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.51 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.35 1.79 0.035 2.12 0.035 2.12 0.26 2.2 0.26 2.2 0.035 2.39 0.035 2.39 0.26 2.47 0.26 2.47 0.035 2.93 0.035 2.93 0.26 3.01 0.26 3.01 0.035 3.205 0.035 3.205 0.255 3.275 0.255 3.275 0.035 3.51 0.035 3.51 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.635 0.035 0.635 0.26 0.715 0.26 0.715 0.035 1.72 0.035 1.72 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 3.51 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.375 1.115 1.375 0.925 1.44 0.925 1.44 0.305 1.375 0.305 1.375 0.085 0.785 0.085 0.785 0.24 0.835 0.24 0.835 0.135 1.04 0.135 1.04 0.255 1.12 0.255 1.12 0.135 1.325 0.135 1.325 0.355 1.39 0.355 1.39 0.875 1.325 0.875 1.325 1.065 1.105 1.065 1.105 0.94 1.055 0.94 1.055 1.065 0.845 1.065 0.845 0.93 0.775 0.93 0.775 1.115 ;
      POLYGON 2.86 1.035 2.86 0.845 2.81 0.845 2.81 0.985 2.59 0.985 2.59 0.925 2.32 0.925 2.32 0.785 2.115 0.785 2.115 0.36 2.59 0.36 2.59 0.17 2.54 0.17 2.54 0.31 2.32 0.31 2.32 0.185 2.27 0.185 2.27 0.31 2.065 0.31 2.065 0.835 2.27 0.835 2.27 0.975 2.54 0.975 2.54 1.035 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 1.25 1.005 1.25 0.825 1.09 0.825 1.09 0.725 0.775 0.725 0.775 0.46 1 0.46 1 0.41 0.725 0.41 0.725 0.775 1.04 0.775 1.04 0.875 1.18 0.875 1.18 1.005 ;
      POLYGON 0.98 1.005 0.98 0.825 0.415 0.825 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.36 1.255 0.36 1.255 0.19 1.175 0.19 1.175 0.31 0.565 0.31 0.565 0.185 0.515 0.185 0.515 0.31 0.365 0.31 0.365 0.425 0.31 0.425 0.31 0.515 0.16 0.515 0.16 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.91 0.875 0.91 1.005 ;
      POLYGON 1.915 0.995 1.915 0.855 1.98 0.855 1.98 0.3 1.915 0.3 1.915 0.16 1.865 0.16 1.865 0.35 1.93 0.35 1.93 0.805 1.865 0.805 1.865 0.995 ;
      POLYGON 1.645 0.97 1.645 0.78 1.575 0.78 1.575 0.35 1.645 0.35 1.645 0.16 1.595 0.16 1.595 0.3 1.525 0.3 1.525 0.83 1.595 0.83 1.595 0.97 ;
      POLYGON 2.725 0.915 2.725 0.775 3.02 0.775 3.02 0.585 3.35 0.585 3.35 0.515 3.02 0.515 3.02 0.31 2.725 0.31 2.725 0.17 2.675 0.17 2.675 0.36 2.97 0.36 2.97 0.725 2.675 0.725 2.675 0.915 ;
      POLYGON 2.6 0.875 2.6 0.675 2.385 0.675 2.385 0.46 2.89 0.46 2.89 0.41 2.335 0.41 2.335 0.515 2.185 0.515 2.185 0.585 2.335 0.585 2.335 0.725 2.54 0.725 2.54 0.825 2.39 0.825 2.39 0.875 ;
      POLYGON 1.05 0.675 1.05 0.53 0.98 0.53 0.98 0.625 0.91 0.625 0.91 0.53 0.84 0.53 0.84 0.675 ;
      RECT 2.44 0.52 2.675 0.6 ;
    LAYER M2 ;
      RECT 1.34 0.825 2.61 0.875 ;
      RECT 0.075 0.825 1.26 0.875 ;
      RECT 0.83 0.625 1.625 0.675 ;
      RECT 1.88 0.525 2.66 0.575 ;
    LAYER VIA1 ;
      RECT 2.43 0.825 2.56 0.875 ;
      RECT 1.39 0.825 1.44 0.875 ;
      RECT 1.08 0.825 1.21 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 1.525 0.625 1.575 0.675 ;
      RECT 0.88 0.625 1.01 0.675 ;
      RECT 2.48 0.525 2.61 0.575 ;
      RECT 1.93 0.525 1.98 0.575 ;
  END
END XOR3_X3M_A12TUL_C35

MACRO XOR3_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.85 0.605 1.85 0.345 1.795 0.345 1.795 0.295 1.645 0.295 1.645 0.085 1.23 0.085 1.23 0.135 1.595 0.135 1.595 0.345 1.745 0.345 1.745 0.395 1.795 0.395 1.795 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.465 0.875 0.465 0.675 0.635 0.675 0.635 0.495 0.58 0.495 0.58 0.625 0.415 0.625 0.415 0.825 0.23 0.825 0.23 0.59 0.175 0.59 0.175 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0287 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.85 0.495 0.85 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0161 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.525 1.01 1.525 0.825 1.31 0.825 1.31 0.445 1.375 0.445 1.375 0.255 1.325 0.255 1.325 0.395 1.255 0.395 1.255 0.875 1.445 0.875 1.445 1.01 ;
    END
    ANTENNADIFFAREA 0.05875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.875 1.72 0.875 1.72 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.31 0.375 0.31 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.715 0.035 1.715 0.245 1.795 0.245 1.795 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.23 0.035 0.23 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.645 1.115 1.645 0.815 1.74 0.815 1.74 0.765 1.595 0.765 1.595 1.065 1.375 1.065 1.375 0.925 1.17 0.925 1.17 0.3 1.255 0.3 1.255 0.22 1.115 0.22 1.115 0.09 1.045 0.09 1.045 0.27 1.12 0.27 1.12 0.925 1.045 0.925 1.045 1.105 1.115 1.105 1.115 0.975 1.325 0.975 1.325 1.115 ;
      POLYGON 0.44 1.105 0.44 0.975 0.565 0.975 0.565 0.755 0.515 0.755 0.515 0.925 0.37 0.925 0.37 1.105 ;
      POLYGON 0.18 1.05 0.18 0.98 0.09 0.98 0.09 0.475 0.415 0.475 0.415 0.155 0.795 0.155 0.795 0.105 0.365 0.105 0.365 0.425 0.16 0.425 0.16 0.22 0.11 0.22 0.11 0.425 0.04 0.425 0.04 1.05 ;
      POLYGON 1.915 1.035 1.915 0.715 1.985 0.715 1.985 0.2 1.85 0.2 1.85 0.28 1.935 0.28 1.935 0.665 1.44 0.665 1.44 0.525 1.39 0.525 1.39 0.715 1.865 0.715 1.865 1.035 ;
      POLYGON 0.72 0.895 0.72 0.875 1.035 0.875 1.035 0.325 0.985 0.325 0.985 0.225 0.485 0.225 0.485 0.275 0.935 0.275 0.935 0.375 0.985 0.375 0.985 0.825 0.63 0.825 0.63 0.895 ;
      POLYGON 0.865 0.775 0.865 0.725 0.75 0.725 0.75 0.375 0.865 0.375 0.865 0.325 0.475 0.325 0.475 0.525 0.31 0.525 0.31 0.715 0.36 0.715 0.36 0.575 0.525 0.575 0.525 0.375 0.7 0.375 0.7 0.775 ;
      POLYGON 1.675 0.445 1.675 0.395 1.51 0.395 1.51 0.255 1.46 0.255 1.46 0.445 ;
  END
END XOR3_X0P5M_A12TUL_C35

MACRO AOI22_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.975 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.445 0.225 0.445 0.085 0.365 0.085 0.365 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.515 0.825 0.515 0.975 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.21 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.635 0.035 0.635 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X0P5M_A12TUL_C35

MACRO NAND2_X0P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.09 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.825 0.245 0.825 0.245 1.09 ;
    END
    ANTENNADIFFAREA 0.03825 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.915 0.1 0.915 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P5B_A12TUL_C35

MACRO XNOR2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.17 0.525 0.22 0.575 ;
        RECT 0.585 0.525 0.635 0.575 ;
      LAYER M1 ;
        RECT 0.565 0.495 0.65 0.675 ;
        RECT 0.16 0.495 0.23 0.775 ;
      LAYER M2 ;
        RECT 0.12 0.525 0.685 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 LAYER M1 ;
    ANTENNAGATEAREA 0.04445 LAYER M2 ;
    ANTENNAGATEAREA 0.04445 LAYER M3 ;
    ANTENNAGATEAREA 0.04445 LAYER M4 ;
    ANTENNAGATEAREA 0.04445 LAYER M5 ;
    ANTENNAGATEAREA 0.04445 LAYER M6 ;
    ANTENNAGATEAREA 0.04445 LAYER M7 ;
    ANTENNAGATEAREA 0.04445 LAYER M8 ;
    ANTENNAGATEAREA 0.04445 LAYER AP ;
    ANTENNAMAXAREACAR 0.9655173 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1231527 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.84 0.395 0.91 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.029575 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.935 0.565 0.775 0.77 0.775 0.77 0.395 0.7 0.395 0.7 0.255 0.65 0.255 0.65 0.445 0.715 0.445 0.715 0.725 0.515 0.725 0.515 0.935 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 1.005 0.235 1.005 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 1 0.235 1 0.185 0.96 0.185 0.96 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.235 0.305 0.235 0.305 0.035 0.89 0.035 0.89 0.235 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.835 1.055 0.835 0.875 1.04 0.875 1.04 0.29 0.835 0.29 0.835 0.23 0.785 0.23 0.785 0.34 0.99 0.34 0.99 0.825 0.785 0.825 0.785 1.005 0.7 1.005 0.7 0.88 0.65 0.88 0.65 1.005 0.43 1.005 0.43 0.885 0.33 0.885 0.33 0.575 0.38 0.575 0.38 0.505 0.28 0.505 0.28 0.935 0.38 0.935 0.38 1.055 ;
      POLYGON 0.16 1.035 0.16 0.845 0.095 0.845 0.095 0.425 0.16 0.425 0.16 0.345 0.43 0.345 0.43 0.135 0.81 0.135 0.81 0.085 0.38 0.085 0.38 0.295 0.16 0.295 0.16 0.235 0.11 0.235 0.11 0.375 0.045 0.375 0.045 0.895 0.11 0.895 0.11 1.035 ;
      POLYGON 0.43 0.815 0.43 0.675 0.5 0.675 0.5 0.445 0.565 0.445 0.565 0.255 0.515 0.255 0.515 0.395 0.35 0.395 0.35 0.445 0.45 0.445 0.45 0.625 0.38 0.625 0.38 0.815 ;
  END
END XNOR2_X1M_A12TUL_C35

MACRO OA21A1OI2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.525 0.235 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.165 0.375 0.165 0.525 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.635 0.505 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.56 0.575 0.56 0.575 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.07 0.7 0.93 0.77 0.93 0.77 0.225 0.575 0.225 0.575 0.09 0.505 0.09 0.505 0.275 0.715 0.275 0.715 0.88 0.65 0.88 0.65 1.07 ;
    END
    ANTENNADIFFAREA 0.037625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.17 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.635 0.035 0.635 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.515 0.875 0.515 1.06 0.565 1.06 0.565 0.825 0.11 0.825 0.11 1.07 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END OA21A1OI2_X0P5M_A12TUL_C35

MACRO NOR2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.31 0.225 0.31 0.095 0.23 0.095 0.23 0.175 0.26 0.175 0.26 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.030125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.175 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.175 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5M_A12TUL_C35

MACRO OAI21_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.565 0.3 0.565 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.635 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01295 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.065 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.065 ;
    END
    ANTENNADIFFAREA 0.03925 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 1 0.505 1 0.505 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END OAI21_X0P5M_A12TUL_C35

MACRO BUF_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.395 0.395 0.395 0.395 0.325 0.175 0.325 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.065 0.43 0.925 0.5 0.925 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.275 0.445 0.275 0.445 0.875 0.38 0.875 0.38 1.065 ;
    END
    ANTENNADIFFAREA 0.03525 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.305 1.165 0.305 0.88 0.235 0.88 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.105 0.17 0.775 0.36 0.775 0.36 0.585 0.31 0.585 0.31 0.725 0.09 0.725 0.09 0.165 0.175 0.165 0.175 0.085 0.04 0.085 0.04 0.775 0.1 0.775 0.1 1.105 ;
  END
END BUF_X0P5M_A12TUL_C35

MACRO AOI21_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.575 0.37 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.3 0.375 0.3 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.425 0.165 0.425 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.495 0.445 0.495 0.445 0.725 0.28 0.725 0.28 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.905 0.635 0.905 0.635 0.225 0.43 0.225 0.43 0.14 0.38 0.14 0.38 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.035375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.21 0.17 0.035 0.5 0.035 0.5 0.17 0.58 0.17 0.58 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.065 0.43 1.065 0.43 0.825 0.11 0.825 0.11 1.07 ;
  END
END AOI21_X0P5M_A12TUL_C35

MACRO BUFH_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.395 0.395 0.395 0.395 0.325 0.175 0.325 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.305 1.165 0.305 0.83 0.235 0.83 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.995 0.16 0.755 0.36 0.755 0.36 0.505 0.31 0.505 0.31 0.705 0.09 0.705 0.09 0.275 0.17 0.275 0.17 0.095 0.1 0.095 0.1 0.225 0.04 0.225 0.04 0.755 0.11 0.755 0.11 0.995 ;
  END
END BUFH_X1M_A12TUL_C35

MACRO OAI31_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI31_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.695 0.665 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.775 0.37 0.565 0.3 0.565 0.3 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.635 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.535 0.64 0.325 0.415 0.325 0.415 0.375 0.57 0.375 0.57 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012075 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.03825 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 1.005 0.64 1.005 0.64 1.165 0.17 1.165 0.17 0.885 0.1 0.885 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.305 0.225 0.305 0.095 0.235 0.095 0.235 0.275 ;
  END
END OAI31_X0P5M_A12TUL_C35

MACRO AOI31_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI31_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013125 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.065 0.7 0.905 0.77 0.905 0.77 0.325 0.575 0.325 0.575 0.09 0.505 0.09 0.505 0.27 0.525 0.27 0.525 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.065 ;
    END
    ANTENNADIFFAREA 0.038125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.64 0.035 0.64 0.175 0.71 0.175 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.055 0.565 0.825 0.245 0.825 0.245 1.055 0.295 1.055 0.295 0.875 0.515 0.875 0.515 1.055 ;
  END
END AOI31_X0P5M_A12TUL_C35

MACRO OAI211_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI211_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.475 0.395 0.475 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.595 0.64 0.395 0.58 0.395 0.58 0.525 0.415 0.525 0.415 0.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.705 0.415 0.705 0.415 0.775 0.615 0.775 0.615 0.825 0.55 0.825 0.55 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 1.11 0.715 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.37 0.925 0.37 1.105 0.44 1.105 0.44 0.975 0.635 0.975 0.635 1.11 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 1.04 0.505 1.04 0.505 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.375 0.43 0.095 0.38 0.095 0.38 0.325 0.17 0.325 0.17 0.09 0.1 0.09 0.1 0.27 0.12 0.27 0.12 0.375 ;
  END
END OAI211_X0P5M_A12TUL_C35

MACRO OAI22_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.44 0.495 0.44 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.775 0.64 0.565 0.57 0.565 0.57 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.06 0.43 0.875 0.77 0.875 0.77 0.325 0.58 0.325 0.58 0.185 0.5 0.185 0.5 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.06 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.925 0.64 0.925 0.64 1.165 0.17 1.165 0.17 0.885 0.1 0.885 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.135 0.65 0.135 0.65 0.22 0.7 0.22 0.7 0.085 0.37 0.085 0.37 0.225 0.16 0.225 0.16 0.11 0.11 0.11 0.11 0.275 ;
  END
END OAI22_X0P5M_A12TUL_C35

MACRO BUF_X1P2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X1P2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.23 0.605 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.02 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.13 0.38 0.13 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.02 ;
    END
    ANTENNADIFFAREA 0.055 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.845 0.235 0.845 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.305 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.045 0.16 0.775 0.495 0.775 0.495 0.585 0.445 0.585 0.445 0.725 0.09 0.725 0.09 0.21 0.18 0.21 0.18 0.14 0.04 0.14 0.04 0.775 0.11 0.775 0.11 1.045 ;
  END
END BUF_X1P2M_A12TUL_C35

MACRO OAI21_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.375 0.725 0.375 0.525 0.295 0.525 0.295 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.655 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.655 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.07675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.58 1.165 0.58 0.93 0.5 0.93 0.5 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OAI21_X1M_A12TUL_C35

MACRO OAI21_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.565 0.3 0.565 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.635 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.58 1.165 0.58 0.93 0.5 0.93 0.5 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OAI21_X0P7M_A12TUL_C35

MACRO OAI21_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.695 0.935 0.625 0.735 0.625 0.735 0.575 0.935 0.575 0.935 0.505 0.685 0.505 0.685 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.095 0.835 0.875 1.04 0.875 1.04 0.325 0.85 0.325 0.85 0.195 0.77 0.195 0.77 0.375 0.985 0.375 0.985 0.825 0.38 0.825 0.38 1.015 0.43 1.015 0.43 0.875 0.785 0.875 0.785 1.095 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 0.375 0.7 0.135 0.91 0.135 0.91 0.27 0.98 0.27 0.98 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.325 0.16 0.325 0.16 0.165 0.11 0.165 0.11 0.375 ;
  END
END OAI21_X1P4M_A12TUL_C35

MACRO OAI22_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.44 0.495 0.44 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.775 0.64 0.565 0.57 0.565 0.57 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.515 0.225 0.515 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.0615 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.925 0.64 0.925 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.275 0.43 0.135 0.64 0.135 0.64 0.27 0.71 0.27 0.71 0.085 0.38 0.085 0.38 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OAI22_X0P7M_A12TUL_C35

MACRO OAI31_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI31_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.695 0.665 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.775 0.37 0.565 0.3 0.565 0.3 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.635 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.565 0.64 0.325 0.415 0.325 0.415 0.375 0.57 0.375 0.57 0.565 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01715 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.985 0.64 0.985 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.305 0.225 0.305 0.095 0.235 0.095 0.235 0.275 ;
  END
END OAI31_X0P7M_A12TUL_C35

MACRO AOI31_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI31_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.325 0.565 0.325 0.565 0.165 0.515 0.165 0.515 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.052625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.64 0.035 0.64 0.2 0.71 0.2 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.015 0.565 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.015 ;
  END
END AOI31_X0P7M_A12TUL_C35

MACRO AO21A1AI2_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.525 0.735 0.525 0.735 0.475 0.8 0.475 0.8 0.425 0.685 0.425 0.685 0.575 0.885 0.575 0.885 0.625 0.715 0.625 0.715 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.205 0.775 1.205 0.705 1.04 0.705 1.04 0.595 1.205 0.595 1.205 0.525 0.985 0.525 0.985 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.19 0.875 1.19 1 1.24 1 1.24 0.875 1.31 0.875 1.31 0.325 1.115 0.325 1.115 0.195 1.045 0.195 1.045 0.375 1.255 0.375 1.255 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.115 1.165 1.115 0.93 1.045 0.93 1.045 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.255 0.845 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.775 0.035 0.775 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.98 1.115 0.98 0.93 0.91 0.93 0.91 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
      POLYGON 0.97 0.375 0.97 0.135 1.18 0.135 1.18 0.27 1.25 0.27 1.25 0.085 0.92 0.085 0.92 0.325 0.7 0.325 0.7 0.175 0.65 0.175 0.65 0.325 0.16 0.325 0.16 0.165 0.11 0.165 0.11 0.375 ;
  END
END AO21A1AI2_X1P4M_A12TUL_C35

MACRO OAI22_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.77 0.875 0.77 0.325 0.575 0.325 0.575 0.195 0.505 0.195 0.505 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.925 0.64 0.925 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.275 0.43 0.135 0.64 0.135 0.64 0.27 0.71 0.27 0.71 0.085 0.38 0.085 0.38 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OAI22_X1M_A12TUL_C35

MACRO AOI21_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.575 0.37 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.3 0.375 0.3 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.425 0.165 0.425 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.495 0.445 0.495 0.445 0.725 0.28 0.725 0.28 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.045 0.565 0.905 0.635 0.905 0.635 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.045 ;
    END
    ANTENNADIFFAREA 0.05 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.5 0.035 0.5 0.17 0.58 0.17 0.58 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.02 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.02 ;
  END
END AOI21_X0P7M_A12TUL_C35

MACRO AOI21_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.575 0.37 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.3 0.375 0.3 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.425 0.165 0.425 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.495 0.445 0.495 0.445 0.725 0.28 0.725 0.28 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.045 0.565 0.905 0.635 0.905 0.635 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.045 ;
    END
    ANTENNADIFFAREA 0.07075 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.5 0.035 0.5 0.17 0.58 0.17 0.58 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.02 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.02 ;
  END
END AOI21_X1M_A12TUL_C35

MACRO OAI31_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI31_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.695 0.665 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.775 0.375 0.525 0.295 0.525 0.295 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.635 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0238 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.07575 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.305 0.225 0.305 0.095 0.235 0.095 0.235 0.275 ;
  END
END OAI31_X1M_A12TUL_C35

MACRO AND3_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND3_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.64 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.64 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.105 0.71 1.005 0.77 1.005 0.77 0.295 0.7 0.295 0.7 0.165 0.65 0.165 0.65 0.355 0.715 0.355 0.715 0.925 0.64 0.925 0.64 1.105 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 1.005 0.235 1.005 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.09 0.16 0.875 0.38 0.875 0.38 1.08 0.43 1.08 0.43 0.875 0.63 0.875 0.63 0.56 0.58 0.56 0.58 0.825 0.08 0.825 0.08 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.03 0.305 0.03 0.875 0.11 0.875 0.11 1.09 ;
  END
END AND3_X0P7M_A12TUL_C35

MACRO OAI211_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI211_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.475 0.395 0.475 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.56 0.175 0.56 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.595 0.64 0.395 0.58 0.395 0.58 0.525 0.415 0.525 0.415 0.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.705 0.415 0.705 0.415 0.775 0.615 0.775 0.615 0.825 0.55 0.825 0.55 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 0.975 0.65 0.975 0.65 1.085 0.7 1.085 0.7 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.061125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 1.035 0.505 1.035 0.505 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.375 0.43 0.175 0.38 0.175 0.38 0.325 0.16 0.325 0.16 0.165 0.11 0.165 0.11 0.375 ;
  END
END OAI211_X0P7M_A12TUL_C35

MACRO AOI22_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.005 0.575 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.505 0.825 0.505 1.005 ;
    END
    ANTENNADIFFAREA 0.0615 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.27 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.635 0.035 0.635 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X0P7M_A12TUL_C35

MACRO OA1B2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA1B2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.235 0.725 0.235 0.525 0.165 0.525 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.805 0.5 0.805 0.5 0.56 0.445 0.56 0.445 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.105 0.71 1.005 0.77 1.005 0.77 0.325 0.565 0.325 0.565 0.13 0.515 0.13 0.515 0.375 0.715 0.375 0.715 0.925 0.64 0.925 0.64 1.105 ;
    END
    ANTENNADIFFAREA 0.0515 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.1 0.16 0.91 0.075 0.91 0.075 0.375 0.415 0.375 0.415 0.475 0.58 0.475 0.58 0.615 0.63 0.615 0.63 0.425 0.465 0.425 0.465 0.325 0.295 0.325 0.295 0.125 0.245 0.125 0.245 0.325 0.025 0.325 0.025 0.96 0.11 0.96 0.11 1.1 ;
  END
END OA1B2_X0P7M_A12TUL_C35

MACRO OA21B_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21B_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.465 0.58 0.465 0.58 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.055 0.7 0.915 0.77 0.915 0.77 0.325 0.565 0.325 0.565 0.13 0.515 0.13 0.515 0.375 0.715 0.375 0.715 0.865 0.65 0.865 0.65 1.055 ;
    END
    ANTENNADIFFAREA 0.0515 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.885 0.37 0.885 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.1 0.16 0.91 0.075 0.91 0.075 0.375 0.415 0.375 0.415 0.515 0.515 0.515 0.515 0.445 0.465 0.445 0.465 0.325 0.295 0.325 0.295 0.125 0.245 0.125 0.245 0.325 0.025 0.325 0.025 0.96 0.11 0.96 0.11 1.1 ;
  END
END OA21B_X0P7M_A12TUL_C35

MACRO OA21A1OI2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.565 0.235 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.165 0.375 0.165 0.565 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.56 0.575 0.56 0.575 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.325 0.565 0.325 0.565 0.165 0.515 0.165 0.515 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.052625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.195 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.64 0.035 0.64 0.195 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.015 0.565 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.515 0.875 0.515 1.015 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OA21A1OI2_X0P7M_A12TUL_C35

MACRO OA21A1OI2_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.625 0.33 0.625 0.33 0.575 0.53 0.575 0.53 0.425 0.31 0.425 0.31 0.475 0.48 0.475 0.48 0.525 0.28 0.525 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.695 0.935 0.505 0.685 0.505 0.685 0.575 0.885 0.575 0.885 0.625 0.685 0.625 0.685 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.205 0.775 1.205 0.705 1.04 0.705 1.04 0.58 1.205 0.58 1.205 0.51 0.985 0.51 0.985 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03605 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.115 1.005 1.115 0.875 1.31 0.875 1.31 0.325 1.24 0.325 1.24 0.185 1.19 0.185 1.19 0.325 0.85 0.325 0.85 0.195 0.77 0.195 0.77 0.375 1.255 0.375 1.255 0.825 1.045 0.825 1.045 1.005 ;
    END
    ANTENNADIFFAREA 0.08825 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 1.115 0.27 1.115 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 1.045 0.035 1.045 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.11 1.25 0.925 1.18 0.925 1.18 1.06 0.97 1.06 0.97 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.11 ;
      POLYGON 0.7 0.375 0.7 0.14 0.91 0.14 0.91 0.27 0.98 0.27 0.98 0.09 0.65 0.09 0.65 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.325 0.16 0.325 0.16 0.165 0.11 0.165 0.11 0.375 ;
  END
END OA21A1OI2_X1P4M_A12TUL_C35

MACRO OAI2XB1_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI2XB1_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.23 0.625 0.23 0.465 0.17 0.465 0.17 0.605 0.145 0.605 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.008225 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.725 0.64 0.725 0.64 0.565 0.57 0.565 0.57 0.725 0.445 0.725 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.775 0.635 0.775 0.425 0.55 0.425 0.55 0.495 0.715 0.495 0.715 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.015 0.7 0.875 0.905 0.875 0.905 0.195 0.845 0.195 0.845 0.095 0.775 0.095 0.775 0.275 0.85 0.275 0.85 0.825 0.65 0.825 0.65 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.44 1.165 0.44 0.835 0.37 0.835 0.37 1.165 0.305 1.165 0.305 1.015 0.235 1.015 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.19 0.17 0.19 0.17 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.175 1.095 0.175 1.015 0.085 1.015 0.085 0.375 0.28 0.375 0.28 0.475 0.445 0.475 0.445 0.615 0.495 0.615 0.495 0.425 0.33 0.425 0.33 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.325 0.035 0.325 0.035 1.095 ;
      POLYGON 0.7 0.375 0.7 0.175 0.65 0.175 0.65 0.325 0.43 0.325 0.43 0.165 0.38 0.165 0.38 0.375 ;
  END
END OAI2XB1_X0P7M_A12TUL_C35

MACRO AOI31_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI31_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.0745 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.015 0.565 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.015 ;
  END
END AOI31_X1M_A12TUL_C35

MACRO INV_X0P6M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P6M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01925 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.065 0.295 0.925 0.365 0.925 0.365 0.26 0.295 0.26 0.295 0.12 0.245 0.12 0.245 0.31 0.31 0.31 0.31 0.875 0.245 0.875 0.245 1.065 ;
    END
    ANTENNADIFFAREA 0.04125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.875 0.1 0.875 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.3 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.3 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P6M_A12TUL_C35

MACRO AOI2XB1_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI2XB1_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.905 0.23 0.675 0.365 0.675 0.365 0.625 0.145 0.625 0.145 0.675 0.175 0.675 0.175 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.635 0.635 0.495 0.665 0.495 0.665 0.425 0.415 0.425 0.415 0.475 0.58 0.475 0.58 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.705 0.55 0.705 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.045 0.835 0.905 0.905 0.905 0.905 0.325 0.7 0.325 0.7 0.13 0.65 0.13 0.65 0.375 0.85 0.375 0.85 0.855 0.785 0.855 0.785 1.045 ;
    END
    ANTENNADIFFAREA 0.05 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 1.015 0.235 1.015 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.315 0.44 0.035 0.775 0.035 0.775 0.195 0.845 0.195 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.175 0.17 0.175 0.17 0.035 0.37 0.035 0.37 0.315 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.18 1.095 0.18 1.025 0.075 1.025 0.075 0.575 0.445 0.575 0.445 0.715 0.495 0.715 0.495 0.525 0.305 0.525 0.305 0.085 0.235 0.085 0.235 0.525 0.025 0.525 0.025 1.095 ;
      POLYGON 0.7 1.015 0.7 0.825 0.38 0.825 0.38 1.015 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1.015 ;
  END
END AOI2XB1_X0P7M_A12TUL_C35

MACRO NAND2_X0P7A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P7A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.095 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.095 ;
    END
    ANTENNADIFFAREA 0.04375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.92 0.1 0.92 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P7A_A12TUL_C35

MACRO BUF_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.395 0.395 0.395 0.395 0.325 0.175 0.325 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0105 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.305 1.165 0.305 0.845 0.235 0.845 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.075 0.16 0.775 0.36 0.775 0.36 0.495 0.31 0.495 0.31 0.725 0.09 0.725 0.09 0.185 0.18 0.185 0.18 0.115 0.04 0.115 0.04 0.775 0.11 0.775 0.11 1.075 ;
  END
END BUF_X1M_A12TUL_C35

MACRO BUF_X9M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X9M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.08085 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.99 0.7 0.88 0.92 0.88 0.92 0.975 0.97 0.975 0.97 0.88 1.19 0.88 1.19 0.975 1.24 0.975 1.24 0.88 1.46 0.88 1.46 0.975 1.51 0.975 1.51 0.88 1.73 0.88 1.73 0.975 1.78 0.975 1.78 0.88 1.865 0.88 1.865 0.32 1.78 0.32 1.78 0.22 1.73 0.22 1.73 0.32 1.51 0.32 1.51 0.225 1.46 0.225 1.46 0.32 1.24 0.32 1.24 0.225 1.19 0.225 1.19 0.32 0.97 0.32 0.97 0.225 0.92 0.225 0.92 0.32 0.7 0.32 0.7 0.21 0.65 0.21 0.65 0.4 1.785 0.4 1.785 0.8 0.65 0.8 0.65 0.99 ;
    END
    ANTENNADIFFAREA 0.437 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.655 1.165 1.655 0.945 1.585 0.945 1.585 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.945 1.045 0.945 1.045 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.355 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.585 0.035 1.585 0.255 1.655 0.255 1.655 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1 0.43 0.875 0.565 0.875 0.565 0.725 0.63 0.725 0.63 0.565 1.65 0.565 1.65 0.605 1.72 0.605 1.72 0.515 0.58 0.515 0.58 0.675 0.515 0.675 0.515 0.825 0.085 0.825 0.085 0.375 0.43 0.375 0.43 0.185 0.38 0.185 0.38 0.325 0.16 0.325 0.16 0.2 0.11 0.2 0.11 0.325 0.035 0.325 0.035 0.875 0.11 0.875 0.11 1 0.16 1 0.16 0.875 0.38 0.875 0.38 1 ;
  END
END BUF_X9M_A12TUL_C35

MACRO BUFH_X6M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X6M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1113 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.015 0.835 0.88 1.055 0.88 1.055 1 1.105 1 1.105 0.88 1.325 0.88 1.325 1 1.375 1 1.375 0.88 1.58 0.88 1.58 0.325 1.375 0.325 1.375 0.205 1.325 0.205 1.325 0.325 1.105 0.325 1.105 0.205 1.055 0.205 1.055 0.325 0.835 0.325 0.835 0.19 0.785 0.19 0.785 0.38 1.525 0.38 1.525 0.825 0.785 0.825 0.785 1.015 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 1.52 1.165 1.52 0.93 1.45 0.93 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.27 1.52 0.27 1.52 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 0.9 0.565 0.775 0.765 0.775 0.765 0.565 1.38 0.565 1.38 0.605 1.45 0.605 1.45 0.515 0.715 0.515 0.715 0.725 0.075 0.725 0.075 0.375 0.565 0.375 0.565 0.185 0.515 0.185 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 0.295 0.9 0.295 0.775 0.515 0.775 0.515 0.9 ;
  END
END BUFH_X6M_A12TUL_C35

MACRO INV_X11M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X11M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.58 0.675 1.58 0.495 1.53 0.495 1.53 0.525 1.175 0.525 1.175 0.425 0.955 0.425 0.955 0.475 1.125 0.475 1.125 0.525 0.635 0.525 0.635 0.425 0.415 0.425 0.415 0.475 0.585 0.475 0.585 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 0.365 0.675 0.365 0.575 0.855 0.575 0.855 0.625 0.685 0.625 0.685 0.675 0.905 0.675 0.905 0.575 1.53 0.575 1.53 0.625 1.36 0.625 1.36 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3542 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.905 0.515 0.905 0.515 0.985 0.565 0.985 0.565 0.905 0.785 0.905 0.785 0.985 0.835 0.985 0.835 0.905 1.055 0.905 1.055 0.985 1.105 0.985 1.105 0.905 1.325 0.905 1.325 0.985 1.375 0.985 1.375 0.905 1.595 0.905 1.595 0.985 1.645 0.985 1.645 0.905 1.73 0.905 1.73 0.28 1.645 0.28 1.645 0.2 1.595 0.2 1.595 0.28 1.375 0.28 1.375 0.2 1.325 0.2 1.325 0.28 1.105 0.28 1.105 0.2 1.055 0.2 1.055 0.28 0.835 0.28 0.835 0.2 0.785 0.2 0.785 0.28 0.565 0.28 0.565 0.2 0.515 0.2 0.515 0.28 0.295 0.28 0.295 0.185 0.245 0.185 0.245 0.375 1.635 0.375 1.635 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
      LAYER M1 ;
        POLYGON 1.755 1.235 1.755 1.165 1.525 1.165 1.525 0.955 1.445 0.955 1.445 1.165 1.255 1.165 1.255 0.955 1.175 0.955 1.175 1.165 0.985 1.165 0.985 0.955 0.905 0.955 0.905 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.755 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.365 0.035 0.365 0.23 0.445 0.23 0.445 0.035 0.635 0.035 0.635 0.23 0.715 0.23 0.715 0.035 0.905 0.035 0.905 0.23 0.985 0.23 0.985 0.035 1.175 0.035 1.175 0.23 1.255 0.23 1.255 0.035 1.445 0.035 1.445 0.23 1.525 0.23 1.525 0.035 1.755 0.035 1.755 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.755 0.065 ;
    END
  END VSS
END INV_X11M_A12TUL_C35

MACRO XNOR3_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.835 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.97 0.425 2.02 0.475 ;
        RECT 2.345 0.425 2.395 0.475 ;
      LAYER M1 ;
        RECT 2.335 0.345 2.405 0.625 ;
        POLYGON 1.99 0.635 1.99 0.495 2.07 0.495 2.07 0.425 1.92 0.425 1.92 0.635 ;
      LAYER M2 ;
        RECT 1.92 0.425 2.445 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01995 LAYER M1 ;
    ANTENNAGATEAREA 0.045675 LAYER M2 ;
    ANTENNAGATEAREA 0.045675 LAYER M3 ;
    ANTENNAGATEAREA 0.045675 LAYER M4 ;
    ANTENNAGATEAREA 0.045675 LAYER M5 ;
    ANTENNAGATEAREA 0.045675 LAYER M6 ;
    ANTENNAGATEAREA 0.045675 LAYER M7 ;
    ANTENNAGATEAREA 0.045675 LAYER M8 ;
    ANTENNAGATEAREA 0.045675 LAYER AP ;
    ANTENNAMAXAREACAR 0.9824563 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1253133 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.505 0.85 0.505 0.85 0.625 0.23 0.625 0.23 0.395 0.175 0.395 0.175 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048125 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.445 0.675 1.445 0.425 1.22 0.425 1.22 0.495 1.39 0.495 1.39 0.625 1.22 0.625 1.22 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04585 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.59 1.015 2.59 0.875 2.795 0.875 2.795 0.325 2.59 0.325 2.59 0.185 2.54 0.185 2.54 0.375 2.74 0.375 2.74 0.825 2.54 0.825 2.54 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
      LAYER M1 ;
        POLYGON 2.835 1.235 2.835 1.165 2.735 1.165 2.735 0.93 2.665 0.93 2.665 1.165 2.47 1.165 2.47 1.03 2.39 1.03 2.39 1.165 1.525 1.165 1.525 1.045 1.445 1.045 1.445 1.165 1.255 1.165 1.255 1.03 1.175 1.03 1.175 1.165 0.575 1.165 0.575 0.845 0.505 0.845 0.505 1.165 0.305 1.165 0.305 0.8 0.235 0.8 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.835 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
      LAYER M1 ;
        POLYGON 2.465 0.275 2.465 0.035 2.665 0.035 2.665 0.27 2.735 0.27 2.735 0.035 2.835 0.035 2.835 -0.035 0 -0.035 0 0.035 0.23 0.035 0.23 0.165 0.31 0.165 0.31 0.035 0.525 0.035 0.525 0.12 0.485 0.12 0.485 0.17 0.595 0.17 0.595 0.035 1.16 0.035 1.16 0.165 1.27 0.165 1.27 0.115 1.23 0.115 1.23 0.035 1.445 0.035 1.445 0.155 1.525 0.155 1.525 0.035 2.395 0.035 2.395 0.275 ;
      LAYER M2 ;
        RECT 0 -0.065 2.835 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.105 1.11 1.105 0.975 1.525 0.975 1.525 0.815 1.575 0.815 1.575 0.325 1.525 0.325 1.525 0.22 0.905 0.22 0.905 0.3 0.985 0.3 0.985 0.27 1.475 0.27 1.475 0.375 1.525 0.375 1.525 0.765 1.475 0.765 1.475 0.925 1.055 0.925 1.055 1.06 0.835 1.06 0.835 0.92 0.785 0.92 0.785 1.11 ;
      POLYGON 1.915 1.065 1.915 0.875 1.71 0.875 1.71 0.27 1.8 0.27 1.8 0.2 1.655 0.2 1.655 0.09 1.585 0.09 1.585 0.27 1.66 0.27 1.66 0.875 1.595 0.875 1.595 1.065 1.645 1.065 1.645 0.925 1.865 0.925 1.865 1.065 ;
      POLYGON 0.16 1.015 0.16 0.825 0.09 0.825 0.09 0.275 0.715 0.275 0.715 0.135 1.08 0.135 1.08 0.085 0.665 0.085 0.665 0.225 0.16 0.225 0.16 0.1 0.11 0.1 0.11 0.225 0.04 0.225 0.04 0.875 0.11 0.875 0.11 1.015 ;
      POLYGON 0.98 1.005 0.98 0.875 1.405 0.875 1.405 0.825 1.105 0.825 1.105 0.37 1.405 0.37 1.405 0.32 1.055 0.32 1.055 0.825 0.91 0.825 0.91 1.005 ;
      POLYGON 2.455 0.975 2.455 0.755 2.52 0.755 2.52 0.575 2.675 0.575 2.675 0.505 2.47 0.505 2.47 0.705 2.405 0.705 2.405 0.925 2.05 0.925 2.05 0.745 1.845 0.745 1.845 0.375 1.925 0.375 1.925 0.195 1.855 0.195 1.855 0.325 1.795 0.325 1.795 0.795 2 0.795 2 0.975 ;
      POLYGON 0.43 0.915 0.43 0.775 0.65 0.775 0.65 0.9 0.7 0.9 0.7 0.775 1.005 0.775 1.005 0.37 0.835 0.37 0.835 0.23 0.785 0.23 0.785 0.325 0.35 0.325 0.35 0.375 0.785 0.375 0.785 0.42 0.955 0.42 0.955 0.725 0.38 0.725 0.38 0.915 ;
      POLYGON 2.33 0.865 2.33 0.685 2.285 0.685 2.285 0.275 2.32 0.275 2.32 0.085 1.755 0.085 1.755 0.135 2.27 0.135 2.27 0.225 2.235 0.225 2.235 0.735 2.26 0.735 2.26 0.865 ;
      POLYGON 2.185 0.865 2.185 0.325 2.06 0.325 2.06 0.195 1.99 0.195 1.99 0.375 2.135 0.375 2.135 0.865 ;
      RECT 0.295 0.505 0.62 0.575 ;
    LAYER M2 ;
      RECT 1.475 0.725 2.235 0.775 ;
      RECT 0.39 0.525 1.155 0.575 ;
    LAYER VIA1 ;
      RECT 2.135 0.725 2.185 0.775 ;
      RECT 1.525 0.725 1.575 0.775 ;
      RECT 1.055 0.525 1.105 0.575 ;
      RECT 0.44 0.525 0.57 0.575 ;
  END
END XNOR3_X2M_A12TUL_C35

MACRO XNOR2_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR2_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.185 0.425 0.235 0.475 ;
        RECT 1.015 0.425 1.145 0.475 ;
      LAYER M1 ;
        POLYGON 1.185 0.625 1.185 0.425 0.975 0.425 0.975 0.625 1.035 0.625 1.035 0.475 1.125 0.475 1.125 0.625 ;
        RECT 0.18 0.375 0.24 0.675 ;
      LAYER M2 ;
        RECT 0.135 0.425 1.195 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 LAYER M1 ;
    ANTENNAGATEAREA 0.0763 LAYER M2 ;
    ANTENNAGATEAREA 0.0763 LAYER M3 ;
    ANTENNAGATEAREA 0.0763 LAYER M4 ;
    ANTENNAGATEAREA 0.0763 LAYER M5 ;
    ANTENNAGATEAREA 0.0763 LAYER M6 ;
    ANTENNAGATEAREA 0.0763 LAYER M7 ;
    ANTENNAGATEAREA 0.0763 LAYER M8 ;
    ANTENNAGATEAREA 0.0763 LAYER AP ;
    ANTENNAMAXAREACAR 0.612245 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2210884 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.805 0.365 0.595 0.53 0.595 0.53 0.525 0.295 0.525 0.295 0.595 0.31 0.595 0.31 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.51 1.105 1.51 0.905 1.58 0.905 1.58 0.295 1.51 0.295 1.51 0.115 0.985 0.115 0.985 0.085 0.905 0.085 0.905 0.165 1.46 0.165 1.46 0.345 1.525 0.345 1.525 0.855 1.46 0.855 1.46 1.055 1.24 1.055 1.24 0.93 1.19 0.93 1.19 1.055 0.985 1.055 0.985 1.025 0.905 1.025 0.905 1.105 ;
    END
    ANTENNADIFFAREA 0.1675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 0.85 1.165 0.85 1.03 0.77 1.03 0.77 1.165 0.575 1.165 0.575 1.045 0.505 1.045 0.505 1.165 0.305 1.165 0.305 0.875 0.235 0.875 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.305 0.305 0.035 0.505 0.035 0.505 0.16 0.575 0.16 0.575 0.035 0.77 0.035 0.77 0.17 0.85 0.17 0.85 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 1.105 0.44 0.975 1.04 0.975 1.04 1 1.12 1 1.12 0.83 1.04 0.83 1.04 0.925 0.55 0.925 0.55 0.725 0.635 0.725 0.635 0.585 0.785 0.585 0.785 0.515 0.635 0.515 0.635 0.425 0.43 0.425 0.43 0.275 1.315 0.275 1.315 0.405 1.385 0.405 1.385 0.225 0.38 0.225 0.38 0.475 0.585 0.475 0.585 0.675 0.5 0.675 0.5 0.925 0.37 0.925 0.37 1.105 ;
      POLYGON 1.375 0.975 1.375 0.725 0.9 0.725 0.9 0.375 1.135 0.375 1.135 0.325 0.62 0.325 0.62 0.375 0.85 0.375 0.85 0.805 0.62 0.805 0.62 0.855 0.9 0.855 0.9 0.775 1.325 0.775 1.325 0.975 ;
      POLYGON 0.16 0.935 0.16 0.745 0.13 0.745 0.13 0.305 0.16 0.305 0.16 0.115 0.11 0.115 0.11 0.255 0.08 0.255 0.08 0.795 0.11 0.795 0.11 0.935 ;
      POLYGON 1.455 0.675 1.455 0.485 1.395 0.485 1.395 0.625 1.305 0.625 1.305 0.485 1.245 0.485 1.245 0.675 ;
    LAYER M2 ;
      RECT 0.04 0.625 1.47 0.675 ;
    LAYER VIA1 ;
      RECT 1.285 0.625 1.415 0.675 ;
      RECT 0.08 0.625 0.13 0.675 ;
  END
END XNOR2_X2M_A12TUL_C35

MACRO XOR2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.805 0.23 0.345 0.43 0.345 0.43 0.135 0.81 0.135 0.81 0.085 0.38 0.085 0.38 0.295 0.175 0.295 0.175 0.405 0.18 0.405 0.18 0.695 0.175 0.695 0.175 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04445 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.845 0.395 0.915 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.029575 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.935 0.565 0.775 0.77 0.775 0.77 0.395 0.7 0.395 0.7 0.255 0.65 0.255 0.65 0.445 0.715 0.445 0.715 0.725 0.515 0.725 0.515 0.935 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 1.005 0.235 1.005 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 1 0.235 1 0.185 0.96 0.185 0.96 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.235 0.305 0.235 0.305 0.035 0.89 0.035 0.89 0.235 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.065 0.16 0.875 0.115 0.875 0.115 0.625 0.13 0.625 0.13 0.475 0.115 0.475 0.115 0.24 0.18 0.24 0.18 0.17 0.065 0.17 0.065 0.925 0.11 0.925 0.11 1.065 ;
      POLYGON 0.835 1.055 0.835 0.875 1.04 0.875 1.04 0.29 0.835 0.29 0.835 0.23 0.785 0.23 0.785 0.34 0.99 0.34 0.99 0.825 0.785 0.825 0.785 1.005 0.7 1.005 0.7 0.88 0.65 0.88 0.65 1.005 0.43 1.005 0.43 0.885 0.33 0.885 0.33 0.575 0.38 0.575 0.38 0.505 0.28 0.505 0.28 0.935 0.38 0.935 0.38 1.055 ;
      POLYGON 0.43 0.815 0.43 0.675 0.5 0.675 0.5 0.445 0.565 0.445 0.565 0.255 0.515 0.255 0.515 0.395 0.35 0.395 0.35 0.445 0.45 0.445 0.45 0.625 0.38 0.625 0.38 0.815 ;
      RECT 0.565 0.495 0.65 0.675 ;
    LAYER M2 ;
      RECT 0.04 0.525 0.685 0.575 ;
    LAYER VIA1 ;
      RECT 0.585 0.525 0.635 0.575 ;
      RECT 0.08 0.525 0.13 0.575 ;
  END
END XOR2_X1M_A12TUL_C35

MACRO XNOR2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.705 0.905 0.425 0.7 0.425 0.7 0.085 0.285 0.085 0.285 0.135 0.65 0.135 0.65 0.475 0.85 0.475 0.85 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0434 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.495 0.175 0.495 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 0.875 0.43 0.735 0.595 0.735 0.595 0.685 0.5 0.685 0.5 0.445 0.565 0.445 0.565 0.23 0.515 0.23 0.515 0.395 0.445 0.395 0.445 0.685 0.38 0.685 0.38 0.875 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.85 1.165 0.85 1.025 0.77 1.025 0.77 1.165 0.17 1.165 0.17 0.895 0.1 0.895 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.355 0.845 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.26 0.17 0.26 0.17 0.035 0.775 0.035 0.775 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 1.105 0.7 0.965 0.97 0.965 0.97 0.825 1.035 0.825 1.035 0.32 0.97 0.32 0.97 0.18 0.92 0.18 0.92 0.37 0.985 0.37 0.985 0.775 0.92 0.775 0.92 0.915 0.65 0.915 0.65 1.055 0.415 1.055 0.415 1.105 ;
      POLYGON 0.565 0.995 0.565 0.855 0.745 0.855 0.745 0.595 0.785 0.595 0.785 0.525 0.695 0.525 0.695 0.805 0.515 0.805 0.515 0.945 0.295 0.945 0.295 0.775 0.085 0.775 0.085 0.375 0.305 0.375 0.305 0.265 0.45 0.265 0.45 0.195 0.235 0.195 0.235 0.325 0.035 0.325 0.035 0.825 0.245 0.825 0.245 0.995 ;
  END
END XNOR2_X0P5M_A12TUL_C35

MACRO BUF_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.014175 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.35 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.095 0.17 0.825 0.33 0.825 0.33 0.745 0.515 0.745 0.515 0.675 0.28 0.675 0.28 0.775 0.09 0.775 0.09 0.27 0.16 0.27 0.16 0.14 0.11 0.14 0.11 0.22 0.04 0.22 0.04 0.825 0.1 0.825 0.1 1.095 ;
  END
END BUF_X1P4M_A12TUL_C35

MACRO AOI22_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.005 0.575 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.505 0.825 0.505 1.005 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.27 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.635 0.035 0.635 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X1M_A12TUL_C35

MACRO NOR2_X0P7A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P7A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.305 0.475 0.305 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.235 0.725 0.235 0.56 0.165 0.56 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.325 0.295 0.325 0.295 0.13 0.245 0.13 0.245 0.375 0.445 0.375 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.0515 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P7A_A12TUL_C35

MACRO NOR2_X1A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X1A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.07325 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.355 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X1A_A12TUL_C35

MACRO XOR2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.105 0.7 0.975 0.835 0.975 0.835 0.805 0.91 0.805 0.91 0.495 0.84 0.495 0.84 0.755 0.785 0.755 0.785 0.925 0.65 0.925 0.65 1.055 0.42 1.055 0.42 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0434 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.495 0.175 0.495 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0245 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 0.875 0.43 0.735 0.595 0.735 0.595 0.685 0.5 0.685 0.5 0.445 0.565 0.445 0.565 0.23 0.515 0.23 0.515 0.395 0.445 0.395 0.445 0.685 0.38 0.685 0.38 0.875 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.85 1.165 0.85 1.03 0.77 1.03 0.77 1.165 0.17 1.165 0.17 0.895 0.1 0.895 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.85 0.33 0.85 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.26 0.17 0.26 0.17 0.035 0.77 0.035 0.77 0.33 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.97 1.065 0.97 0.925 1.035 0.925 1.035 0.385 0.97 0.385 0.97 0.23 0.92 0.23 0.92 0.385 0.7 0.385 0.7 0.085 0.285 0.085 0.285 0.135 0.65 0.135 0.65 0.435 0.985 0.435 0.985 0.875 0.92 0.875 0.92 1.065 ;
      POLYGON 0.565 0.995 0.565 0.855 0.715 0.855 0.715 0.595 0.785 0.595 0.785 0.525 0.665 0.525 0.665 0.805 0.515 0.805 0.515 0.945 0.295 0.945 0.295 0.775 0.085 0.775 0.085 0.375 0.305 0.375 0.305 0.265 0.45 0.265 0.45 0.195 0.235 0.195 0.235 0.325 0.035 0.325 0.035 0.825 0.245 0.825 0.245 0.995 ;
  END
END XOR2_X0P5M_A12TUL_C35

MACRO XOR3_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 4.59 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 2.075 0.525 2.125 0.575 ;
        RECT 3.31 0.525 3.44 0.575 ;
      LAYER M1 ;
        RECT 2.06 0.43 2.14 0.645 ;
        POLYGON 3.48 0.655 3.48 0.525 3.27 0.525 3.27 0.655 3.34 0.655 3.34 0.575 3.41 0.575 3.41 0.655 ;
      LAYER M2 ;
        RECT 2.025 0.525 3.49 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 LAYER M1 ;
    ANTENNAGATEAREA 0.08995 LAYER M2 ;
    ANTENNAGATEAREA 0.08995 LAYER M3 ;
    ANTENNAGATEAREA 0.08995 LAYER M4 ;
    ANTENNAGATEAREA 0.08995 LAYER M5 ;
    ANTENNAGATEAREA 0.08995 LAYER M6 ;
    ANTENNAGATEAREA 0.08995 LAYER M7 ;
    ANTENNAGATEAREA 0.08995 LAYER M8 ;
    ANTENNAGATEAREA 0.08995 LAYER AP ;
    ANTENNAMAXAREACAR 0.5341615 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2018634 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.295 0.625 1.425 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 1.455 0.685 1.455 0.505 1.385 0.505 1.385 0.615 1.32 0.615 1.32 0.505 1.25 0.505 1.25 0.685 ;
        POLYGON 1.99 0.685 1.99 0.525 1.92 0.525 1.92 0.615 1.855 0.615 1.855 0.505 1.785 0.505 1.785 0.685 ;
      LAYER M2 ;
        RECT 1.245 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04165 LAYER M1 ;
    ANTENNAGATEAREA 0.09135 LAYER M2 ;
    ANTENNAGATEAREA 0.09135 LAYER M3 ;
    ANTENNAGATEAREA 0.09135 LAYER M4 ;
    ANTENNAGATEAREA 0.09135 LAYER M5 ;
    ANTENNAGATEAREA 0.09135 LAYER M6 ;
    ANTENNAGATEAREA 0.09135 LAYER M7 ;
    ANTENNAGATEAREA 0.09135 LAYER M8 ;
    ANTENNAGATEAREA 0.09135 LAYER AP ;
    ANTENNAMAXAREACAR 0.6806723 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1560625 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.675 0.665 0.625 0.465 0.625 0.465 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.067725 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 1.015 4.075 0.875 4.295 0.875 4.295 1.005 4.345 1.005 4.345 0.875 4.55 0.875 4.55 0.325 4.345 0.325 4.345 0.19 4.295 0.19 4.295 0.325 4.075 0.325 4.075 0.185 4.025 0.185 4.025 0.375 4.495 0.375 4.495 0.825 4.025 0.825 4.025 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
        RECT 3.485 1.175 3.535 1.225 ;
        RECT 3.62 1.175 3.67 1.225 ;
        RECT 3.755 1.175 3.805 1.225 ;
        RECT 3.89 1.175 3.94 1.225 ;
        RECT 4.025 1.175 4.075 1.225 ;
        RECT 4.16 1.175 4.21 1.225 ;
        RECT 4.295 1.175 4.345 1.225 ;
        RECT 4.43 1.175 4.48 1.225 ;
      LAYER M1 ;
        POLYGON 4.59 1.235 4.59 1.165 4.49 1.165 4.49 0.93 4.42 0.93 4.42 1.165 4.22 1.165 4.22 0.945 4.15 0.945 4.15 1.165 3.95 1.165 3.95 0.845 3.88 0.845 3.88 1.165 3.145 1.165 3.145 1.03 3.065 1.03 3.065 1.165 2.87 1.165 2.87 0.775 2.8 0.775 2.8 1.165 2.6 1.165 2.6 0.93 2.53 0.93 2.53 1.165 2.33 1.165 2.33 0.93 2.26 0.93 2.26 1.165 2.06 1.165 2.06 0.795 1.99 0.795 1.99 1.165 1.79 1.165 1.79 0.875 1.72 0.875 1.72 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 4.59 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
        RECT 3.485 -0.025 3.535 0.025 ;
        RECT 3.62 -0.025 3.67 0.025 ;
        RECT 3.755 -0.025 3.805 0.025 ;
        RECT 3.89 -0.025 3.94 0.025 ;
        RECT 4.025 -0.025 4.075 0.025 ;
        RECT 4.16 -0.025 4.21 0.025 ;
        RECT 4.295 -0.025 4.345 0.025 ;
        RECT 4.43 -0.025 4.48 0.025 ;
      LAYER M1 ;
        POLYGON 2.06 0.36 2.06 0.035 2.26 0.035 2.26 0.27 2.33 0.27 2.33 0.035 2.53 0.035 2.53 0.335 2.6 0.335 2.6 0.035 2.8 0.035 2.8 0.27 2.87 0.27 2.87 0.035 3.07 0.035 3.07 0.27 3.14 0.27 3.14 0.035 3.88 0.035 3.88 0.35 3.95 0.35 3.95 0.035 4.15 0.035 4.15 0.255 4.22 0.255 4.22 0.035 4.42 0.035 4.42 0.27 4.49 0.27 4.49 0.035 4.59 0.035 4.59 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.72 0.035 1.72 0.305 1.79 0.305 1.79 0.035 1.99 0.035 1.99 0.36 ;
      LAYER M2 ;
        RECT 0 -0.065 4.59 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.51 1.115 1.51 0.925 1.575 0.925 1.575 0.385 1.51 0.385 1.51 0.26 1.46 0.26 1.46 0.385 1.24 0.385 1.24 0.185 0.91 0.185 0.91 0.365 0.98 0.365 0.98 0.235 1.19 0.235 1.19 0.435 1.525 0.435 1.525 0.875 1.46 0.875 1.46 1.065 1.24 1.065 1.24 0.94 1.19 0.94 1.19 1.065 0.97 1.065 0.97 0.965 0.92 0.965 0.92 1.115 ;
      POLYGON 3.67 1.105 3.67 0.915 3.62 0.915 3.62 1.055 3.265 1.055 3.265 0.925 2.995 0.925 2.995 0.655 2.79 0.655 2.79 0.375 3.41 0.375 3.41 0.195 3.34 0.195 3.34 0.325 2.995 0.325 2.995 0.2 2.945 0.2 2.945 0.325 2.74 0.325 2.74 0.705 2.945 0.705 2.945 0.975 3.215 0.975 3.215 1.105 ;
      POLYGON 0.835 1.02 0.835 0.895 1.04 0.895 1.04 1.005 1.12 1.005 1.12 0.845 0.415 0.845 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.375 0.835 0.375 0.835 0.135 1.325 0.135 1.325 0.325 1.375 0.325 1.375 0.085 0.785 0.085 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.365 0.325 0.365 0.425 0.31 0.425 0.31 0.515 0.16 0.515 0.16 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.895 0.515 0.895 0.515 1.02 0.565 1.02 0.565 0.895 0.785 0.895 0.785 1.02 ;
      POLYGON 2.455 1.015 2.455 0.875 2.675 0.875 2.675 0.405 2.455 0.405 2.455 0.265 2.405 0.265 2.405 0.455 2.625 0.455 2.625 0.825 2.405 0.825 2.405 1.015 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 3.41 1.005 3.41 0.825 3.115 0.825 3.115 0.475 3.67 0.475 3.67 0.23 3.62 0.23 3.62 0.425 3.065 0.425 3.065 0.515 2.86 0.515 2.86 0.585 3.065 0.585 3.065 0.875 3.34 0.875 3.34 1.005 ;
      POLYGON 1.385 1.005 1.385 0.825 1.225 0.825 1.225 0.745 0.9 0.745 0.9 0.475 1.12 0.475 1.12 0.29 1.04 0.29 1.04 0.425 0.85 0.425 0.85 0.795 1.175 0.795 1.175 0.875 1.315 0.875 1.315 1.005 ;
      POLYGON 1.915 1 1.915 0.745 1.71 0.745 1.71 0.425 1.915 0.425 1.915 0.165 1.865 0.165 1.865 0.375 1.66 0.375 1.66 0.795 1.865 0.795 1.865 1 ;
      POLYGON 3.805 0.9 3.805 0.775 3.875 0.775 3.875 0.575 4.34 0.575 4.34 0.595 4.43 0.595 4.43 0.525 3.875 0.525 3.875 0.42 3.805 0.42 3.805 0.085 3.205 0.085 3.205 0.27 3.275 0.27 3.275 0.135 3.485 0.135 3.485 0.26 3.535 0.26 3.535 0.135 3.755 0.135 3.755 0.47 3.825 0.47 3.825 0.725 3.185 0.725 3.185 0.775 3.485 0.775 3.485 0.9 3.535 0.9 3.535 0.775 3.755 0.775 3.755 0.9 ;
      POLYGON 2.185 0.89 2.185 0.75 2.25 0.75 2.25 0.325 2.185 0.325 2.185 0.185 2.135 0.185 2.135 0.375 2.2 0.375 2.2 0.7 2.135 0.7 2.135 0.89 ;
      POLYGON 2.355 0.875 2.355 0.595 2.54 0.595 2.54 0.525 2.305 0.525 2.305 0.805 2.245 0.805 2.245 0.875 ;
      POLYGON 1.19 0.685 1.19 0.525 0.97 0.525 0.97 0.685 1.05 0.685 1.05 0.595 1.11 0.595 1.11 0.685 ;
      POLYGON 3.75 0.675 3.75 0.545 3.68 0.545 3.68 0.625 3.61 0.625 3.61 0.545 3.54 0.545 3.54 0.675 ;
    LAYER M2 ;
      RECT 2.455 0.825 3.285 0.875 ;
      RECT 1.475 0.825 2.375 0.875 ;
      RECT 0.075 0.825 1.395 0.875 ;
      RECT 2.15 0.625 3.76 0.675 ;
      RECT 0.965 0.525 1.76 0.575 ;
    LAYER VIA1 ;
      RECT 3.105 0.825 3.235 0.875 ;
      RECT 2.505 0.825 2.635 0.875 ;
      RECT 2.275 0.825 2.325 0.875 ;
      RECT 1.525 0.825 1.575 0.875 ;
      RECT 1.215 0.825 1.345 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 3.58 0.625 3.71 0.675 ;
      RECT 2.2 0.625 2.25 0.675 ;
      RECT 1.66 0.525 1.71 0.575 ;
      RECT 1.015 0.525 1.145 0.575 ;
  END
END XOR3_X4M_A12TUL_C35

MACRO XOR2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.19 0.425 0.24 0.475 ;
        RECT 0.485 0.425 0.615 0.475 ;
      LAYER M1 ;
        POLYGON 0.5 0.6 0.5 0.475 0.71 0.475 0.71 0.54 0.78 0.54 0.78 0.425 0.435 0.425 0.435 0.6 ;
        RECT 0.18 0.375 0.25 0.695 ;
      LAYER M2 ;
        RECT 0.14 0.425 0.665 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02835 LAYER M1 ;
    ANTENNAGATEAREA 0.0574 LAYER M2 ;
    ANTENNAGATEAREA 0.0574 LAYER M3 ;
    ANTENNAGATEAREA 0.0574 LAYER M4 ;
    ANTENNAGATEAREA 0.0574 LAYER M5 ;
    ANTENNAGATEAREA 0.0574 LAYER M6 ;
    ANTENNAGATEAREA 0.0574 LAYER M7 ;
    ANTENNAGATEAREA 0.0574 LAYER M8 ;
    ANTENNAGATEAREA 0.0574 LAYER AP ;
    ANTENNAMAXAREACAR 1.055556 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.229277 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.465 0.85 0.465 0.85 0.605 0.715 0.605 0.715 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0308 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.005 0.575 0.875 1.04 0.875 1.04 0.325 0.72 0.325 0.72 0.3 0.63 0.3 0.63 0.375 0.985 0.375 0.985 0.825 0.505 0.825 0.505 1.005 ;
    END
    ANTENNADIFFAREA 0.079 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.91 0.035 0.91 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.845 1.11 0.845 0.93 0.775 0.93 0.775 1.06 0.71 1.06 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.36 0.825 0.36 0.375 0.565 0.375 0.565 0.25 0.85 0.25 0.85 0.09 0.77 0.09 0.77 0.2 0.515 0.2 0.515 0.325 0.31 0.325 0.31 0.875 0.38 0.875 0.38 1.11 ;
      POLYGON 0.16 0.98 0.16 0.79 0.13 0.79 0.13 0.305 0.16 0.305 0.16 0.115 0.11 0.115 0.11 0.25 0.08 0.25 0.08 0.84 0.11 0.84 0.11 0.98 ;
      POLYGON 0.65 0.775 0.65 0.53 0.57 0.53 0.57 0.725 0.43 0.725 0.43 0.775 ;
      POLYGON 0.44 0.27 0.44 0.15 0.595 0.15 0.595 0.09 0.37 0.09 0.37 0.27 ;
    LAYER M2 ;
      RECT 0.04 0.725 0.655 0.775 ;
    LAYER VIA1 ;
      RECT 0.475 0.725 0.605 0.775 ;
      RECT 0.08 0.725 0.13 0.775 ;
  END
END XOR2_X0P7M_A12TUL_C35

MACRO NAND2_X2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0602 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0602 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.131 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X2B_A12TUL_C35

MACRO NAND2_X1A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.06175 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X1A_A12TUL_C35

MACRO OR2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OR2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.565 0.17 0.565 0.17 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.017675 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.305 0.475 0.305 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.017675 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.045 0.565 0.905 0.635 0.905 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.045 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.835 0.37 0.835 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.025 0.16 0.835 0.075 0.835 0.075 0.375 0.445 0.375 0.445 0.595 0.495 0.595 0.495 0.325 0.295 0.325 0.295 0.12 0.245 0.12 0.245 0.325 0.025 0.325 0.025 0.885 0.11 0.885 0.11 1.025 ;
  END
END OR2_X1M_A12TUL_C35

MACRO CGENI_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN CGENI_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.495 0.58 0.495 0.58 0.625 0.24 0.625 0.24 0.525 0.16 0.525 0.16 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.575 0.53 0.505 0.365 0.505 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.005 0.71 0.875 0.905 0.875 0.905 0.325 0.71 0.325 0.71 0.195 0.64 0.195 0.64 0.375 0.85 0.375 0.85 0.825 0.64 0.825 0.64 1.005 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END CON
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.845 1.115 0.845 0.93 0.775 0.93 0.775 1.065 0.565 1.065 0.565 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.115 ;
      POLYGON 0.565 0.375 0.565 0.135 0.775 0.135 0.775 0.27 0.845 0.27 0.845 0.085 0.515 0.085 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 ;
  END
END CGENI_X1M_A12TUL_C35

MACRO XNOR3_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.51 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.795 0.625 1.845 0.675 ;
        RECT 2.785 0.625 2.835 0.675 ;
      LAYER M1 ;
        POLYGON 2.91 0.675 2.91 0.605 2.815 0.605 2.815 0.515 2.735 0.515 2.735 0.675 ;
        RECT 1.785 0.42 1.855 0.71 ;
      LAYER M2 ;
        RECT 1.745 0.625 2.885 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 LAYER M1 ;
    ANTENNAGATEAREA 0.05495 LAYER M2 ;
    ANTENNAGATEAREA 0.05495 LAYER M3 ;
    ANTENNAGATEAREA 0.05495 LAYER M4 ;
    ANTENNAGATEAREA 0.05495 LAYER M5 ;
    ANTENNAGATEAREA 0.05495 LAYER M6 ;
    ANTENNAGATEAREA 0.05495 LAYER M7 ;
    ANTENNAGATEAREA 0.05495 LAYER M8 ;
    ANTENNAGATEAREA 0.05495 LAYER AP ;
    ANTENNAMAXAREACAR 0.8923078 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1098901 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.88 0.525 1.01 0.575 ;
        RECT 1.66 0.525 1.71 0.575 ;
      LAYER M1 ;
        POLYGON 1.05 0.65 1.05 0.525 0.84 0.525 0.84 0.65 0.91 0.65 0.91 0.575 0.98 0.575 0.98 0.65 ;
        RECT 1.65 0.42 1.72 0.71 ;
      LAYER M2 ;
        RECT 0.83 0.525 1.76 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0308 LAYER M1 ;
    ANTENNAGATEAREA 0.0924 LAYER M2 ;
    ANTENNAGATEAREA 0.0924 LAYER M3 ;
    ANTENNAGATEAREA 0.0924 LAYER M4 ;
    ANTENNAGATEAREA 0.0924 LAYER M5 ;
    ANTENNAGATEAREA 0.0924 LAYER M6 ;
    ANTENNAGATEAREA 0.0924 LAYER M7 ;
    ANTENNAGATEAREA 0.0924 LAYER M8 ;
    ANTENNAGATEAREA 0.0924 LAYER AP ;
    ANTENNAMAXAREACAR 0.659091 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.211039 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.465 0.625 0.465 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05775 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 3.13 1.015 3.13 0.875 3.35 0.875 3.35 1 3.4 1 3.4 0.875 3.47 0.875 3.47 0.325 3.4 0.325 3.4 0.2 3.35 0.2 3.35 0.325 3.13 0.325 3.13 0.185 3.08 0.185 3.08 0.375 3.415 0.375 3.415 0.825 3.08 0.825 3.08 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
      LAYER M1 ;
        POLYGON 3.51 1.235 3.51 1.165 3.275 1.165 3.275 0.945 3.205 0.945 3.205 1.165 3.005 1.165 3.005 0.845 2.935 0.845 2.935 1.165 2.47 1.165 2.47 1.03 2.39 1.03 2.39 1.165 2.195 1.165 2.195 0.905 2.125 0.905 2.125 1.165 1.79 1.165 1.79 0.78 1.72 0.78 1.72 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.925 0.1 0.925 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.51 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.35 1.79 0.035 2.12 0.035 2.12 0.26 2.2 0.26 2.2 0.035 2.39 0.035 2.39 0.26 2.47 0.26 2.47 0.035 2.93 0.035 2.93 0.26 3.01 0.26 3.01 0.035 3.205 0.035 3.205 0.255 3.275 0.255 3.275 0.035 3.51 0.035 3.51 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.635 0.035 0.635 0.26 0.715 0.26 0.715 0.035 1.72 0.035 1.72 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 3.51 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.375 1.115 1.375 0.925 1.445 0.925 1.445 0.325 1.375 0.325 1.375 0.09 0.785 0.09 0.785 0.24 0.835 0.24 0.835 0.14 1.04 0.14 1.04 0.26 1.12 0.26 1.12 0.14 1.325 0.14 1.325 0.375 1.395 0.375 1.395 0.875 1.325 0.875 1.325 1.065 1.105 1.065 1.105 0.94 1.055 0.94 1.055 1.065 0.845 1.065 0.845 0.93 0.775 0.93 0.775 1.115 ;
      POLYGON 2.86 1.035 2.86 0.845 2.81 0.845 2.81 0.985 2.59 0.985 2.59 0.925 2.32 0.925 2.32 0.785 2.115 0.785 2.115 0.36 2.59 0.36 2.59 0.17 2.54 0.17 2.54 0.31 2.32 0.31 2.32 0.185 2.27 0.185 2.27 0.31 2.065 0.31 2.065 0.835 2.27 0.835 2.27 0.975 2.54 0.975 2.54 1.035 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 1.25 1.005 1.25 0.825 1.09 0.825 1.09 0.725 0.775 0.725 0.775 0.465 1 0.465 1 0.415 0.725 0.415 0.725 0.775 1.04 0.775 1.04 0.875 1.18 0.875 1.18 1.005 ;
      POLYGON 0.98 1.005 0.98 0.825 0.415 0.825 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.36 1.255 0.36 1.255 0.2 1.175 0.2 1.175 0.31 0.565 0.31 0.565 0.185 0.515 0.185 0.515 0.31 0.365 0.31 0.365 0.425 0.31 0.425 0.31 0.515 0.16 0.515 0.16 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.91 0.875 0.91 1.005 ;
      POLYGON 1.915 0.995 1.915 0.855 1.98 0.855 1.98 0.3 1.915 0.3 1.915 0.16 1.865 0.16 1.865 0.35 1.93 0.35 1.93 0.805 1.865 0.805 1.865 0.995 ;
      POLYGON 1.645 0.97 1.645 0.78 1.575 0.78 1.575 0.35 1.645 0.35 1.645 0.16 1.595 0.16 1.595 0.3 1.525 0.3 1.525 0.83 1.595 0.83 1.595 0.97 ;
      POLYGON 2.725 0.915 2.725 0.775 3.02 0.775 3.02 0.585 3.35 0.585 3.35 0.515 3.02 0.515 3.02 0.31 2.725 0.31 2.725 0.17 2.675 0.17 2.675 0.36 2.97 0.36 2.97 0.725 2.675 0.725 2.675 0.915 ;
      POLYGON 2.6 0.875 2.6 0.665 2.385 0.665 2.385 0.46 2.89 0.46 2.89 0.41 2.335 0.41 2.335 0.515 2.185 0.515 2.185 0.585 2.335 0.585 2.335 0.715 2.54 0.715 2.54 0.825 2.39 0.825 2.39 0.875 ;
      POLYGON 1.32 0.675 1.32 0.52 1.25 0.52 1.25 0.625 1.18 0.625 1.18 0.52 1.11 0.52 1.11 0.675 ;
      RECT 2.44 0.52 2.675 0.6 ;
    LAYER M2 ;
      RECT 1.345 0.825 2.61 0.875 ;
      RECT 0.075 0.825 1.26 0.875 ;
      RECT 1.1 0.625 1.625 0.675 ;
      RECT 1.88 0.525 2.66 0.575 ;
    LAYER VIA1 ;
      RECT 2.43 0.825 2.56 0.875 ;
      RECT 1.395 0.825 1.445 0.875 ;
      RECT 1.08 0.825 1.21 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 1.525 0.625 1.575 0.675 ;
      RECT 1.15 0.625 1.28 0.675 ;
      RECT 2.48 0.525 2.61 0.575 ;
      RECT 1.93 0.525 1.98 0.575 ;
  END
END XNOR3_X3M_A12TUL_C35

MACRO AO21A1AI2_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.525 0.735 0.525 0.735 0.475 0.8 0.475 0.8 0.425 0.685 0.425 0.685 0.575 0.885 0.575 0.885 0.625 0.715 0.625 0.715 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.205 0.775 1.205 0.705 1.04 0.705 1.04 0.595 1.205 0.595 1.205 0.525 0.985 0.525 0.985 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04655 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.19 0.875 1.19 1 1.24 1 1.24 0.875 1.31 0.875 1.31 0.325 1.115 0.325 1.115 0.195 1.045 0.195 1.045 0.375 1.255 0.375 1.255 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.13025 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.115 1.165 1.115 0.93 1.045 0.93 1.045 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.255 0.845 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.775 0.035 0.775 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.98 1.115 0.98 0.93 0.91 0.93 0.91 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
      POLYGON 0.97 0.375 0.97 0.135 1.18 0.135 1.18 0.27 1.25 0.27 1.25 0.085 0.92 0.085 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END AO21A1AI2_X2M_A12TUL_C35

MACRO MXIT2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN MXIT2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.495 0.31 0.495 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.705 0.77 0.495 0.8 0.495 0.8 0.425 0.685 0.425 0.685 0.495 0.71 0.495 0.71 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.55 0.63 0.55 0.63 0.44 0.58 0.44 0.58 0.495 0.445 0.495 0.445 0.725 0.23 0.725 0.23 0.565 0.175 0.565 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03395 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 0.975 0.715 0.975 0.715 0.875 0.905 0.875 0.905 0.325 0.71 0.325 0.71 0.225 0.575 0.225 0.575 0.095 0.505 0.095 0.505 0.275 0.66 0.275 0.66 0.375 0.85 0.375 0.85 0.825 0.665 0.825 0.665 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.059 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.05 0.16 0.875 0.61 0.875 0.61 0.735 0.65 0.735 0.65 0.665 0.56 0.665 0.56 0.825 0.085 0.825 0.085 0.375 0.445 0.375 0.445 0.435 0.495 0.435 0.495 0.325 0.16 0.325 0.16 0.15 0.11 0.15 0.11 0.325 0.035 0.325 0.035 0.875 0.11 0.875 0.11 1.05 ;
  END
END MXIT2_X0P5M_A12TUL_C35

MACRO OAI21_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.845 0.325 0.845 0.195 0.775 0.195 0.775 0.375 0.985 0.375 0.985 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 0.375 0.7 0.135 0.91 0.135 0.91 0.27 0.98 0.27 0.98 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OAI21_X2M_A12TUL_C35

MACRO INV_X2P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X2P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.080325 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.133875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X2P5M_A12TUL_C35

MACRO OAI2XB1_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI2XB1_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.23 0.625 0.23 0.465 0.175 0.465 0.175 0.605 0.145 0.605 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0105 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.725 0.645 0.725 0.645 0.525 0.565 0.525 0.565 0.725 0.445 0.725 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.775 0.645 0.775 0.425 0.55 0.425 0.55 0.475 0.715 0.475 0.715 0.645 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.015 0.7 0.875 0.905 0.875 0.905 0.295 0.835 0.295 0.835 0.155 0.785 0.155 0.785 0.345 0.85 0.345 0.85 0.825 0.65 0.825 0.65 1.015 ;
    END
    ANTENNADIFFAREA 0.07675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.44 1.165 0.44 0.835 0.37 0.835 0.37 1.165 0.305 1.165 0.305 1 0.235 1 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.19 0.17 0.19 0.17 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.175 1.06 0.175 0.98 0.085 0.98 0.085 0.375 0.28 0.375 0.28 0.575 0.425 0.575 0.425 0.595 0.515 0.595 0.515 0.525 0.33 0.525 0.33 0.325 0.295 0.325 0.295 0.1 0.245 0.1 0.245 0.325 0.035 0.325 0.035 1.06 ;
      POLYGON 0.7 0.375 0.7 0.185 0.65 0.185 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 ;
  END
END OAI2XB1_X1M_A12TUL_C35

MACRO OA21A1OI2_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.625 0.33 0.625 0.33 0.575 0.53 0.575 0.53 0.425 0.31 0.425 0.31 0.475 0.48 0.475 0.48 0.525 0.28 0.525 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.525 0.735 0.525 0.735 0.475 0.8 0.475 0.8 0.425 0.685 0.425 0.685 0.575 0.885 0.575 0.885 0.625 0.715 0.625 0.715 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.205 0.775 1.205 0.705 1.04 0.705 1.04 0.58 1.205 0.58 1.205 0.51 0.985 0.51 0.985 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05005 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.115 1.005 1.115 0.875 1.31 0.875 1.31 0.325 1.24 0.325 1.24 0.2 1.19 0.2 1.19 0.325 0.845 0.325 0.845 0.195 0.775 0.195 0.775 0.375 1.255 0.375 1.255 0.825 1.045 0.825 1.045 1.005 ;
    END
    ANTENNADIFFAREA 0.12275 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 1.115 0.27 1.115 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 1.045 0.035 1.045 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.11 1.25 0.925 1.18 0.925 1.18 1.06 0.97 1.06 0.97 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.11 ;
      POLYGON 0.7 0.375 0.7 0.14 0.91 0.14 0.91 0.27 0.98 0.27 0.98 0.09 0.65 0.09 0.65 0.325 0.43 0.325 0.43 0.195 0.38 0.195 0.38 0.325 0.16 0.325 0.16 0.18 0.11 0.18 0.11 0.375 ;
  END
END OA21A1OI2_X2M_A12TUL_C35

MACRO NOR2_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.575 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.505 0.28 0.505 0.28 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03605 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03605 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.77 0.875 0.77 0.225 0.565 0.225 0.565 0.125 0.515 0.125 0.515 0.225 0.295 0.225 0.295 0.125 0.245 0.125 0.245 0.275 0.715 0.275 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.067 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.2 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.635 0.035 0.635 0.17 0.715 0.17 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.2 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NOR2_X1P4M_A12TUL_C35

MACRO NAND2B_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2B_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.55 0.175 0.55 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.11 0.44 0.975 0.635 0.975 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.27 0.58 0.27 0.58 0.925 0.37 0.925 0.37 1.11 ;
    END
    ANTENNADIFFAREA 0.04075 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.58 1.165 0.58 1.03 0.5 1.03 0.5 1.165 0.305 1.165 0.305 0.995 0.235 0.995 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.175 1.1 0.175 1.02 0.075 1.02 0.075 0.375 0.445 0.375 0.445 0.57 0.495 0.57 0.495 0.325 0.175 0.325 0.175 0.085 0.095 0.085 0.095 0.325 0.025 0.325 0.025 1.1 ;
  END
END NAND2B_X0P7M_A12TUL_C35

MACRO AOI211_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI211_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.225 0.715 0.225 0.715 0.09 0.635 0.09 0.635 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.715 0.275 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.05925 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.505 0.035 0.505 0.165 0.575 0.165 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.02 0.43 0.825 0.11 0.825 0.11 1.02 0.16 1.02 0.16 0.875 0.38 0.875 0.38 1.02 ;
  END
END AOI211_X0P7M_A12TUL_C35

MACRO AND3_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND3_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.64 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.64 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.105 0.71 1.005 0.77 1.005 0.77 0.215 0.71 0.215 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.64 0.925 0.64 1.105 ;
    END
    ANTENNADIFFAREA 0.034875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 1.02 0.235 1.02 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.105 0.17 0.875 0.37 0.875 0.37 1.095 0.44 1.095 0.44 0.875 0.63 0.875 0.63 0.665 0.58 0.665 0.58 0.825 0.08 0.825 0.08 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.03 0.305 0.03 0.875 0.1 0.875 0.1 1.105 ;
  END
END AND3_X0P5M_A12TUL_C35

MACRO OAI21B_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21B_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.635 0.645 0.425 0.415 0.425 0.415 0.475 0.575 0.475 0.575 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.485 0.715 0.485 0.715 0.705 0.55 0.705 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.575 0.365 0.525 0.23 0.525 0.23 0.295 0.175 0.295 0.175 0.505 0.145 0.505 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.905 0.875 0.905 0.325 0.43 0.325 0.43 0.165 0.38 0.165 0.38 0.375 0.85 0.375 0.85 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.44 1.165 0.44 0.92 0.37 0.92 0.37 1.165 0.305 1.165 0.305 1.01 0.235 1.01 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.18 0.305 0.035 0.64 0.035 0.64 0.165 0.71 0.165 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.105 0.16 0.775 0.495 0.775 0.495 0.57 0.445 0.57 0.445 0.725 0.085 0.725 0.085 0.175 0.175 0.175 0.175 0.095 0.035 0.095 0.035 0.775 0.11 0.775 0.11 1.105 ;
      POLYGON 0.845 0.275 0.845 0.095 0.775 0.095 0.775 0.225 0.575 0.225 0.575 0.095 0.505 0.095 0.505 0.275 ;
  END
END OAI21B_X0P7M_A12TUL_C35

MACRO AOI2XB1_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI2XB1_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.905 0.23 0.675 0.365 0.675 0.365 0.625 0.145 0.625 0.145 0.675 0.175 0.675 0.175 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.635 0.635 0.495 0.665 0.495 0.665 0.425 0.415 0.425 0.415 0.475 0.58 0.475 0.58 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.705 0.55 0.705 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.07 0.835 0.905 0.905 0.905 0.905 0.325 0.7 0.325 0.7 0.14 0.65 0.14 0.65 0.375 0.85 0.375 0.85 0.855 0.785 0.855 0.785 1.07 ;
    END
    ANTENNADIFFAREA 0.035375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 1.015 0.235 1.015 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.21 0.44 0.035 0.775 0.035 0.775 0.175 0.845 0.175 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.175 0.17 0.175 0.17 0.035 0.37 0.035 0.37 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.18 1.095 0.18 1.025 0.075 1.025 0.075 0.575 0.445 0.575 0.445 0.715 0.495 0.715 0.495 0.525 0.305 0.525 0.305 0.085 0.235 0.085 0.235 0.525 0.025 0.525 0.025 1.095 ;
      POLYGON 0.43 1.07 0.43 0.875 0.65 0.875 0.65 1.055 0.7 1.055 0.7 0.825 0.38 0.825 0.38 1.07 ;
  END
END AOI2XB1_X0P5M_A12TUL_C35

MACRO NOR2B_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2B_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.235 0.725 0.235 0.525 0.165 0.525 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.008925 ;
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.635 0.375 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.325 0.43 0.325 0.43 0.11 0.38 0.11 0.38 0.375 0.58 0.375 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.06025 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.305 1.165 0.305 0.93 0.235 0.93 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.09 0.16 0.875 0.495 0.875 0.495 0.505 0.445 0.505 0.445 0.825 0.075 0.825 0.075 0.175 0.18 0.175 0.18 0.105 0.025 0.105 0.025 0.875 0.11 0.875 0.11 1.09 ;
  END
END NOR2B_X1M_A12TUL_C35

MACRO AND2_X0P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND2_X0P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007525 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.325 0.145 0.325 0.145 0.375 0.31 0.375 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007525 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.09 0.5 0.09 0.5 0.17 0.58 0.17 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.027 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0.17 1.165 0.17 1.025 0.1 1.025 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.17 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.305 1.105 0.305 0.875 0.495 0.875 0.495 0.225 0.175 0.225 0.175 0.085 0.095 0.085 0.095 0.165 0.125 0.165 0.125 0.275 0.445 0.275 0.445 0.825 0.255 0.825 0.255 1.015 0.235 1.015 0.235 1.105 ;
  END
END AND2_X0P5B_A12TUL_C35

MACRO OAI2XB1_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI2XB1_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.23 0.625 0.23 0.465 0.17 0.465 0.17 0.605 0.145 0.605 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.007875 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.725 0.64 0.725 0.64 0.565 0.57 0.565 0.57 0.725 0.445 0.725 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.635 0.77 0.425 0.55 0.425 0.55 0.495 0.715 0.495 0.715 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.07 0.7 0.875 0.905 0.875 0.905 0.195 0.845 0.195 0.845 0.09 0.775 0.09 0.775 0.27 0.85 0.27 0.85 0.825 0.65 0.825 0.65 1.07 ;
    END
    ANTENNADIFFAREA 0.03875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 1.005 0.775 1.005 0.775 1.165 0.44 1.165 0.44 0.885 0.37 0.885 0.37 1.165 0.305 1.165 0.305 1.02 0.235 1.02 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.175 1.1 0.175 1.02 0.085 1.02 0.085 0.375 0.28 0.375 0.28 0.475 0.445 0.475 0.445 0.615 0.495 0.615 0.495 0.425 0.33 0.425 0.33 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.325 0.035 0.325 0.035 1.1 ;
      POLYGON 0.7 0.375 0.7 0.095 0.65 0.095 0.65 0.325 0.44 0.325 0.44 0.09 0.37 0.09 0.37 0.27 0.39 0.27 0.39 0.375 ;
  END
END OAI2XB1_X0P5M_A12TUL_C35

MACRO AO21B_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.62 0.375 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.62 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.705 0.635 0.705 0.635 0.495 0.58 0.495 0.58 0.705 0.445 0.705 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.095 0.64 0.095 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.07575 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.835 0.37 0.835 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.095 0.295 0.825 0.075 0.825 0.075 0.355 0.445 0.355 0.445 0.605 0.495 0.605 0.495 0.305 0.16 0.305 0.16 0.16 0.11 0.16 0.11 0.305 0.025 0.305 0.025 0.875 0.245 0.875 0.245 1.095 ;
  END
END AO21B_X1M_A12TUL_C35

MACRO XNOR2_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR2_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.7 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.55 0.525 1.68 0.575 ;
        RECT 2.36 0.525 2.49 0.575 ;
      LAYER M1 ;
        RECT 1.375 0.525 1.73 0.595 ;
        POLYGON 2.52 0.705 2.52 0.515 2.33 0.515 2.33 0.705 2.385 0.705 2.385 0.585 2.47 0.585 2.47 0.705 ;
      LAYER M2 ;
        RECT 1.5 0.525 2.54 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 LAYER M1 ;
    ANTENNAGATEAREA 0.13545 LAYER M2 ;
    ANTENNAGATEAREA 0.13545 LAYER M3 ;
    ANTENNAGATEAREA 0.13545 LAYER M4 ;
    ANTENNAGATEAREA 0.13545 LAYER M5 ;
    ANTENNAGATEAREA 0.13545 LAYER M6 ;
    ANTENNAGATEAREA 0.13545 LAYER M7 ;
    ANTENNAGATEAREA 0.13545 LAYER M8 ;
    ANTENNAGATEAREA 0.13545 LAYER AP ;
    ANTENNAMAXAREACAR 0.560606 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1406928 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 1.205 0.575 1.205 0.425 0.955 0.425 0.955 0.475 1.155 0.475 1.155 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.05 1 2.05 0.875 2.255 0.875 2.255 0.325 2.05 0.325 2.05 0.2 2 0.2 2 0.325 1.78 0.325 1.78 0.185 1.45 0.185 1.45 0.365 1.52 0.365 1.52 0.235 1.73 0.235 1.73 0.375 2.2 0.375 2.2 0.825 1.915 0.825 1.915 0.725 1.43 0.725 1.43 0.775 1.865 0.775 1.865 0.875 2 0.875 2 1 ;
    END
    ANTENNADIFFAREA 0.255 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
      LAYER M1 ;
        POLYGON 2.7 1.235 2.7 1.165 2.6 1.165 2.6 0.905 2.53 0.905 2.53 1.165 2.33 1.165 2.33 0.925 2.26 0.925 2.26 1.165 1.255 1.165 1.255 1.03 1.175 1.03 1.175 1.165 0.98 1.165 0.98 0.845 0.91 0.845 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.7 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.175 0.035 1.175 0.17 1.255 0.17 1.255 0.035 2.26 0.035 2.26 0.275 2.33 0.275 2.33 0.035 2.53 0.035 2.53 0.325 2.6 0.325 2.6 0.035 2.7 0.035 2.7 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.7 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 2.195 1.115 2.195 0.93 2.125 0.93 2.125 1.065 1.915 1.065 1.915 0.925 1.78 0.925 1.78 0.825 1.305 0.825 1.305 0.475 1.655 0.475 1.655 0.285 1.585 0.285 1.585 0.425 1.375 0.425 1.375 0.345 1.325 0.345 1.325 0.425 1.255 0.425 1.255 0.875 1.73 0.875 1.73 0.975 1.865 0.975 1.865 1.115 ;
      POLYGON 1.655 1.105 1.655 0.925 1.105 0.925 1.105 0.725 0.63 0.725 0.63 0.475 0.835 0.475 0.835 0.375 1.105 0.375 1.105 0.275 1.375 0.275 1.375 0.135 1.865 0.135 1.865 0.26 1.915 0.26 1.915 0.135 2.125 0.135 2.125 0.275 2.195 0.275 2.195 0.085 1.325 0.085 1.325 0.225 1.105 0.225 1.105 0.185 1.055 0.185 1.055 0.325 0.835 0.325 0.835 0.275 0.785 0.275 0.785 0.425 0.58 0.425 0.58 0.525 0.15 0.525 0.15 0.575 0.58 0.575 0.58 0.775 0.785 0.775 0.785 0.9 0.835 0.9 0.835 0.775 1.055 0.775 1.055 0.975 1.325 0.975 1.325 1.1 1.375 1.1 1.375 0.975 1.585 0.975 1.585 1.105 ;
      POLYGON 0.565 1.015 0.565 0.825 0.09 0.825 0.09 0.375 0.565 0.375 0.565 0.185 0.515 0.185 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1 0.295 1 0.295 0.875 0.515 0.875 0.515 1.015 ;
      POLYGON 2.455 0.975 2.455 0.835 2.62 0.835 2.62 0.395 2.455 0.395 2.455 0.195 2.405 0.195 2.405 0.445 2.57 0.445 2.57 0.785 2.405 0.785 2.405 0.975 ;
      POLYGON 2.12 0.675 2.12 0.565 2.07 0.565 2.07 0.625 1.985 0.625 1.985 0.565 1.935 0.565 1.935 0.625 1.85 0.625 1.85 0.565 1.8 0.565 1.8 0.675 ;
    LAYER M2 ;
      RECT 0.335 0.825 1.49 0.875 ;
      RECT 1.89 0.625 2.66 0.675 ;
    LAYER VIA1 ;
      RECT 1.31 0.825 1.44 0.875 ;
      RECT 0.385 0.825 0.515 0.875 ;
      RECT 2.57 0.625 2.62 0.675 ;
      RECT 1.94 0.625 2.07 0.675 ;
  END
END XNOR2_X4M_A12TUL_C35

MACRO NAND2_X1P4A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1P4A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.425 0.28 0.425 0.28 0.495 0.445 0.495 0.445 0.605 0.28 0.605 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.095 0.565 0.875 0.77 0.875 0.77 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.095 0.295 1.095 0.295 0.875 0.515 0.875 0.515 1.095 ;
    END
    ANTENNADIFFAREA 0.073 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.94 0.37 0.94 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X1P4A_A12TUL_C35

MACRO NAND3_X0P5A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND3_X0P5A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.37 0.825 0.37 0.625 0.3 0.625 0.3 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.775 0.235 0.575 0.365 0.575 0.365 0.525 0.145 0.525 0.145 0.575 0.165 0.575 0.165 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.095 0.565 0.975 0.635 0.975 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.27 0.58 0.27 0.58 0.925 0.245 0.925 0.245 1.085 0.295 1.085 0.295 0.975 0.515 0.975 0.515 1.095 ;
    END
    ANTENNADIFFAREA 0.041125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 1.035 0.37 1.035 0.37 1.165 0.17 1.165 0.17 1.01 0.1 1.01 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END NAND3_X0P5A_A12TUL_C35

MACRO NOR3_X0P5A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR3_X0P5A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.875 0.5 0.595 0.445 0.595 0.445 0.825 0.28 0.825 0.28 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013475 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013475 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013475 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.225 0.575 0.225 0.575 0.1 0.505 0.1 0.505 0.225 0.295 0.225 0.295 0.1 0.245 0.1 0.245 0.275 0.58 0.275 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.041875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.185 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.185 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END NOR3_X0P5A_A12TUL_C35

MACRO OA21B_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21B_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.465 0.58 0.465 0.58 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.055 0.7 0.915 0.77 0.915 0.77 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.715 0.375 0.715 0.865 0.65 0.865 0.65 1.055 ;
    END
    ANTENNADIFFAREA 0.07325 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.22 0.17 0.22 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.04 0.16 0.835 0.075 0.835 0.075 0.375 0.415 0.375 0.415 0.515 0.515 0.515 0.515 0.445 0.465 0.445 0.465 0.325 0.305 0.325 0.305 0.09 0.235 0.09 0.235 0.325 0.025 0.325 0.025 0.885 0.11 0.885 0.11 1.04 ;
  END
END OA21B_X1M_A12TUL_C35

MACRO AOI21_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03605 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.125 0.785 0.125 0.785 0.325 0.43 0.325 0.43 0.14 0.38 0.14 0.38 0.375 0.985 0.375 0.985 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.077 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.315 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.2 0.98 0.2 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.315 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.98 1.115 0.98 0.93 0.91 0.93 0.91 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
  END
END AOI21_X1P4M_A12TUL_C35

MACRO MX2_X2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN MX2_X2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.775 0.8 0.725 0.635 0.725 0.635 0.675 0.8 0.675 0.8 0.625 0.58 0.625 0.58 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.235 0.725 0.235 0.565 0.165 0.565 0.165 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.615 0.365 0.475 0.5 0.475 0.5 0.325 0.28 0.325 0.28 0.375 0.43 0.375 0.43 0.425 0.31 0.425 0.31 0.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.033425 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.105 1.015 1.105 0.875 1.325 0.875 1.325 1 1.375 1 1.375 0.875 1.58 0.875 1.58 0.325 1.375 0.325 1.375 0.225 1.25 0.225 1.25 0.095 1.18 0.095 1.18 0.275 1.325 0.275 1.325 0.375 1.525 0.375 1.525 0.825 1.055 0.825 1.055 1.015 ;
    END
    ANTENNADIFFAREA 0.131 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 1.52 1.165 1.52 0.93 1.45 0.93 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.925 0.37 0.925 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 1.52 0.27 1.52 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.45 0.035 1.45 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.065 0.565 0.825 0.52 0.825 0.52 0.575 0.84 0.575 0.84 0.595 0.925 0.595 0.925 0.525 0.6 0.525 0.6 0.115 0.5 0.115 0.5 0.195 0.55 0.195 0.55 0.525 0.47 0.525 0.47 0.875 0.515 0.875 0.515 1.065 ;
      POLYGON 0.835 1.025 0.835 0.885 0.97 0.885 0.97 0.735 1.165 0.735 1.165 0.615 1.325 0.615 1.325 0.545 1.165 0.545 1.165 0.325 0.7 0.325 0.7 0.175 0.65 0.175 0.65 0.375 1.115 0.375 1.115 0.685 0.92 0.685 0.92 0.835 0.785 0.835 0.785 1.025 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.495 0.26 0.495 0.26 0.425 0.16 0.425 0.16 0.18 0.11 0.18 0.11 0.425 0.04 0.425 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 1.45 0.605 1.45 0.425 1.235 0.425 1.235 0.475 1.395 0.475 1.395 0.605 ;
      POLYGON 1.04 0.595 1.04 0.425 0.82 0.425 0.82 0.475 0.99 0.475 0.99 0.595 ;
    LAYER M2 ;
      RECT 0.04 0.425 1.455 0.475 ;
    LAYER VIA1 ;
      RECT 1.275 0.425 1.405 0.475 ;
      RECT 0.86 0.425 0.99 0.475 ;
      RECT 0.09 0.425 0.22 0.475 ;
  END
END MX2_X2B_A12TUL_C35

MACRO ADDF_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN ADDF_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.295 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.595 0.625 0.725 0.675 ;
        RECT 1.255 0.625 1.305 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 0.765 0.675 0.765 0.505 0.715 0.505 0.715 0.625 0.36 0.625 0.36 0.505 0.31 0.505 0.31 0.675 ;
        POLYGON 1.335 0.675 1.335 0.605 1.315 0.605 1.315 0.415 1.245 0.415 1.245 0.605 1.225 0.605 1.225 0.675 ;
        POLYGON 1.855 0.725 1.855 0.675 2 0.675 2 0.625 1.855 0.625 1.855 0.535 1.785 0.535 1.785 0.725 ;
      LAYER M2 ;
        RECT 0.545 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.10465 LAYER M2 ;
    ANTENNAGATEAREA 0.10465 LAYER M3 ;
    ANTENNAGATEAREA 0.10465 LAYER M4 ;
    ANTENNAGATEAREA 0.10465 LAYER M5 ;
    ANTENNAGATEAREA 0.10465 LAYER M6 ;
    ANTENNAGATEAREA 0.10465 LAYER M7 ;
    ANTENNAGATEAREA 0.10465 LAYER M8 ;
    ANTENNAGATEAREA 0.10465 LAYER AP ;
    ANTENNAMAXAREACAR 1.304762 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.475 0.425 0.605 0.475 ;
        RECT 1.425 0.425 1.555 0.475 ;
        RECT 1.825 0.425 1.955 0.475 ;
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.425 0.435 0.425 0.435 0.575 0.505 0.575 0.505 0.475 0.575 0.475 0.575 0.575 ;
        POLYGON 1.995 0.575 1.995 0.425 1.785 0.425 1.785 0.475 1.925 0.475 1.925 0.575 ;
        POLYGON 1.455 0.605 1.455 0.475 1.595 0.475 1.595 0.425 1.385 0.425 1.385 0.605 ;
      LAYER M2 ;
        RECT 0.425 0.425 2.005 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.10465 LAYER M2 ;
    ANTENNAGATEAREA 0.10465 LAYER M3 ;
    ANTENNAGATEAREA 0.10465 LAYER M4 ;
    ANTENNAGATEAREA 0.10465 LAYER M5 ;
    ANTENNAGATEAREA 0.10465 LAYER M6 ;
    ANTENNAGATEAREA 0.10465 LAYER M7 ;
    ANTENNAGATEAREA 0.10465 LAYER M8 ;
    ANTENNAGATEAREA 0.10465 LAYER AP ;
    ANTENNAMAXAREACAR 1.111111 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.85 0.525 0.9 0.575 ;
        RECT 1.11 0.525 1.16 0.575 ;
        RECT 1.665 0.525 1.715 0.575 ;
      LAYER M1 ;
        RECT 0.84 0.42 0.91 0.675 ;
        RECT 1.1 0.415 1.17 0.685 ;
        RECT 1.665 0.445 1.715 0.755 ;
      LAYER M2 ;
        RECT 0.8 0.525 1.765 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.07245 LAYER M2 ;
    ANTENNAGATEAREA 0.07245 LAYER M3 ;
    ANTENNAGATEAREA 0.07245 LAYER M4 ;
    ANTENNAGATEAREA 0.07245 LAYER M5 ;
    ANTENNAGATEAREA 0.07245 LAYER M6 ;
    ANTENNAGATEAREA 0.07245 LAYER M7 ;
    ANTENNAGATEAREA 0.07245 LAYER M8 ;
    ANTENNAGATEAREA 0.07245 LAYER AP ;
    ANTENNAMAXAREACAR 0.984127 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1587302 LAYER VIA1 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.17 1.105 0.17 0.925 0.095 0.925 0.095 0.27 0.17 0.27 0.17 0.09 0.1 0.09 0.1 0.195 0.04 0.195 0.04 1.005 0.1 1.005 0.1 1.105 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.195 1.105 2.195 1.005 2.255 1.005 2.255 0.195 2.195 0.195 2.195 0.09 2.125 0.09 2.125 0.27 2.2 0.27 2.2 0.925 2.125 0.925 2.125 1.105 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
      LAYER M1 ;
        POLYGON 2.295 1.235 2.295 1.165 2.06 1.165 2.06 0.905 1.99 0.905 1.99 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.855 1.045 0.855 1.045 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.855 0.235 0.855 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.295 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.375 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 1.045 0.035 1.045 0.27 1.115 0.27 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.295 0.035 2.295 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.295 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.97 1.065 0.97 0.875 0.92 0.875 0.92 1.015 0.7 1.015 0.7 0.845 0.38 0.845 0.38 1.035 0.43 1.035 0.43 0.895 0.65 0.895 0.65 1.065 ;
      POLYGON 1.645 1.045 1.645 0.905 1.845 0.905 1.845 0.835 2.12 0.835 2.12 0.325 1.645 0.325 1.645 0.165 1.595 0.165 1.595 0.375 2.07 0.375 2.07 0.785 1.795 0.785 1.795 0.855 1.595 0.855 1.595 1.045 ;
      POLYGON 1.51 1.035 1.51 0.845 1.19 0.845 1.19 1.035 1.24 1.035 1.24 0.895 1.46 0.895 1.46 1.035 ;
      POLYGON 0.835 0.91 0.835 0.785 1.58 0.785 1.58 0.605 1.53 0.605 1.53 0.735 1.035 0.735 1.035 0.32 0.845 0.32 0.845 0.19 0.775 0.19 0.775 0.37 0.985 0.37 0.985 0.735 0.225 0.735 0.225 0.505 0.175 0.505 0.175 0.785 0.785 0.785 0.785 0.91 ;
      POLYGON 0.7 0.375 0.7 0.135 0.91 0.135 0.91 0.27 0.98 0.27 0.98 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 ;
      POLYGON 1.51 0.355 1.51 0.165 1.46 0.165 1.46 0.305 1.24 0.305 1.24 0.165 1.19 0.165 1.19 0.355 ;
  END
END ADDF_X1M_A12TUL_C35

MACRO BUF_X13M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X13M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.7 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1162 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 0.96 0.835 0.885 1.055 0.885 1.055 0.945 1.105 0.945 1.105 0.885 1.325 0.885 1.325 0.945 1.375 0.945 1.375 0.885 1.595 0.885 1.595 0.945 1.645 0.945 1.645 0.885 1.865 0.885 1.865 0.945 1.915 0.945 1.915 0.885 2.135 0.885 2.135 0.945 2.185 0.945 2.185 0.885 2.405 0.885 2.405 0.945 2.455 0.945 2.455 0.885 2.59 0.885 2.59 0.285 2.54 0.285 2.54 0.315 2.455 0.315 2.455 0.25 2.405 0.25 2.405 0.315 2.185 0.315 2.185 0.25 2.135 0.25 2.135 0.315 1.915 0.315 1.915 0.25 1.865 0.25 1.865 0.315 1.645 0.315 1.645 0.25 1.595 0.25 1.595 0.315 1.375 0.315 1.375 0.25 1.325 0.25 1.325 0.315 1.105 0.315 1.105 0.25 1.055 0.25 1.055 0.315 0.835 0.315 0.835 0.24 0.785 0.24 0.785 0.43 2.47 0.43 2.47 0.77 0.785 0.77 0.785 0.96 ;
    END
    ANTENNADIFFAREA 0.713 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
      LAYER M1 ;
        POLYGON 2.7 1.235 2.7 1.165 2.33 1.165 2.33 0.945 2.26 0.945 2.26 1.165 2.06 1.165 2.06 0.945 1.99 0.945 1.99 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.7 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 1.72 0.035 1.72 0.255 1.79 0.255 1.79 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.26 0.035 2.26 0.255 2.33 0.255 2.33 0.035 2.7 0.035 2.7 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.7 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1 0.565 0.875 0.7 0.875 0.7 0.71 0.77 0.71 0.77 0.565 2.325 0.565 2.325 0.605 2.395 0.605 2.395 0.515 0.72 0.515 0.72 0.66 0.65 0.66 0.65 0.825 0.085 0.825 0.085 0.375 0.565 0.375 0.565 0.185 0.515 0.185 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.035 0.325 0.035 0.875 0.245 0.875 0.245 1 0.295 1 0.295 0.875 0.515 0.875 0.515 1 ;
  END
END BUF_X13M_A12TUL_C35

MACRO NOR2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.56 0.175 0.56 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018025 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.445 1.11 0.445 1.005 0.5 1.005 0.5 0.225 0.295 0.225 0.295 0.125 0.245 0.125 0.245 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.11 ;
    END
    ANTENNADIFFAREA 0.0425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.195 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P7M_A12TUL_C35

MACRO XOR2_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.7 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.94 0.625 2.07 0.675 ;
        RECT 2.36 0.625 2.49 0.675 ;
      LAYER M1 ;
        POLYGON 2.12 0.675 2.12 0.565 2.07 0.565 2.07 0.625 1.985 0.625 1.985 0.565 1.935 0.565 1.935 0.625 1.85 0.625 1.85 0.565 1.8 0.565 1.8 0.675 ;
        POLYGON 2.52 0.685 2.52 0.495 2.47 0.495 2.47 0.615 2.385 0.615 2.385 0.495 2.33 0.495 2.33 0.685 ;
      LAYER M2 ;
        RECT 1.89 0.625 2.54 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 LAYER M1 ;
    ANTENNAGATEAREA 0.13545 LAYER M2 ;
    ANTENNAGATEAREA 0.13545 LAYER M3 ;
    ANTENNAGATEAREA 0.13545 LAYER M4 ;
    ANTENNAGATEAREA 0.13545 LAYER M5 ;
    ANTENNAGATEAREA 0.13545 LAYER M6 ;
    ANTENNAGATEAREA 0.13545 LAYER M7 ;
    ANTENNAGATEAREA 0.13545 LAYER M8 ;
    ANTENNAGATEAREA 0.13545 LAYER AP ;
    ANTENNAMAXAREACAR 0.560606 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1406928 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 1.205 0.575 1.205 0.425 0.985 0.425 0.985 0.475 1.155 0.475 1.155 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.05 1 2.05 0.875 2.255 0.875 2.255 0.325 2.05 0.325 2.05 0.2 2 0.2 2 0.325 1.78 0.325 1.78 0.185 1.45 0.185 1.45 0.365 1.52 0.365 1.52 0.235 1.73 0.235 1.73 0.375 2.2 0.375 2.2 0.825 1.915 0.825 1.915 0.725 1.43 0.725 1.43 0.775 1.865 0.775 1.865 0.875 2 0.875 2 1 ;
    END
    ANTENNADIFFAREA 0.255 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
      LAYER M1 ;
        POLYGON 2.7 1.235 2.7 1.165 2.6 1.165 2.6 0.875 2.53 0.875 2.53 1.165 2.33 1.165 2.33 0.925 2.26 0.925 2.26 1.165 1.255 1.165 1.255 1.03 1.175 1.03 1.175 1.165 0.98 1.165 0.98 0.845 0.91 0.845 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.7 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.18 1.25 0.18 1.25 0.035 2.26 0.035 2.26 0.275 2.33 0.275 2.33 0.035 2.53 0.035 2.53 0.305 2.6 0.305 2.6 0.035 2.7 0.035 2.7 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.7 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 2.195 1.115 2.195 0.93 2.125 0.93 2.125 1.065 1.915 1.065 1.915 0.925 1.78 0.925 1.78 0.825 1.31 0.825 1.31 0.475 1.655 0.475 1.655 0.29 1.585 0.29 1.585 0.425 1.375 0.425 1.375 0.36 1.325 0.36 1.325 0.425 1.26 0.425 1.26 0.875 1.73 0.875 1.73 0.975 1.865 0.975 1.865 1.115 ;
      POLYGON 1.655 1.105 1.655 0.925 1.105 0.925 1.105 0.725 0.63 0.725 0.63 0.475 0.835 0.475 0.835 0.375 1.105 0.375 1.105 0.3 1.375 0.3 1.375 0.135 1.865 0.135 1.865 0.26 1.915 0.26 1.915 0.135 2.125 0.135 2.125 0.275 2.195 0.275 2.195 0.085 1.325 0.085 1.325 0.25 1.105 0.25 1.105 0.185 1.055 0.185 1.055 0.325 0.835 0.325 0.835 0.275 0.785 0.275 0.785 0.425 0.58 0.425 0.58 0.525 0.15 0.525 0.15 0.575 0.58 0.575 0.58 0.775 0.785 0.775 0.785 0.9 0.835 0.9 0.835 0.775 1.055 0.775 1.055 0.975 1.325 0.975 1.325 1.1 1.375 1.1 1.375 0.975 1.585 0.975 1.585 1.105 ;
      POLYGON 0.565 1.015 0.565 0.825 0.09 0.825 0.09 0.375 0.565 0.375 0.565 0.185 0.515 0.185 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1 0.295 1 0.295 0.875 0.515 0.875 0.515 1.015 ;
      POLYGON 2.455 0.965 2.455 0.805 2.62 0.805 2.62 0.375 2.455 0.375 2.455 0.195 2.405 0.195 2.405 0.425 2.57 0.425 2.57 0.755 2.405 0.755 2.405 0.965 ;
      RECT 1.375 0.525 1.73 0.595 ;
    LAYER M2 ;
      RECT 0.335 0.825 1.49 0.875 ;
      RECT 1.5 0.525 2.66 0.575 ;
    LAYER VIA1 ;
      RECT 1.31 0.825 1.44 0.875 ;
      RECT 0.385 0.825 0.515 0.875 ;
      RECT 2.57 0.525 2.62 0.575 ;
      RECT 1.55 0.525 1.68 0.575 ;
  END
END XOR2_X4M_A12TUL_C35

MACRO AOI22BB_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22BB_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.625 0.77 0.625 0.77 0.445 0.715 0.445 0.715 0.625 0.58 0.625 0.58 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.585 0.905 0.325 0.685 0.325 0.685 0.375 0.85 0.375 0.85 0.585 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END B0N
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.705 0.23 0.705 0.23 0.545 0.175 0.545 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0133 ;
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.965 0.565 0.775 1.04 0.775 1.04 0.225 0.71 0.225 0.71 0.095 0.64 0.095 0.64 0.275 0.985 0.275 0.985 0.725 0.515 0.725 0.515 0.965 ;
    END
    ANTENNADIFFAREA 0.054125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.17 1.165 0.17 0.915 0.1 0.915 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.27 0.575 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.37 0.035 0.37 0.195 0.44 0.195 0.44 0.035 0.505 0.035 0.505 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.105 0.43 0.96 0.465 0.96 0.465 0.555 0.65 0.555 0.65 0.485 0.465 0.485 0.465 0.305 0.295 0.305 0.295 0.125 0.245 0.125 0.245 0.355 0.415 0.355 0.415 0.91 0.38 0.91 0.38 1.105 ;
      POLYGON 0.97 1.015 0.97 0.825 0.65 0.825 0.65 1.015 0.7 1.015 0.7 0.875 0.92 0.875 0.92 1.015 ;
  END
END AOI22BB_X0P7M_A12TUL_C35

MACRO OAI211_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI211_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.475 0.395 0.475 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.555 0.175 0.555 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.595 0.64 0.395 0.58 0.395 0.58 0.525 0.415 0.525 0.415 0.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021875 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.705 0.415 0.705 0.415 0.775 0.615 0.775 0.615 0.825 0.55 0.825 0.55 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021875 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.11 0.71 0.975 0.77 0.975 0.77 0.275 0.7 0.275 0.7 0.135 0.65 0.135 0.65 0.325 0.715 0.325 0.715 0.925 0.37 0.925 0.37 1.105 0.44 1.105 0.44 0.975 0.64 0.975 0.64 1.11 ;
    END
    ANTENNADIFFAREA 0.08675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 1.035 0.505 1.035 0.505 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.375 0.43 0.18 0.38 0.18 0.38 0.325 0.16 0.325 0.16 0.18 0.11 0.18 0.11 0.375 ;
  END
END OAI211_X1M_A12TUL_C35

MACRO AOI2XB1_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI2XB1_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.905 0.23 0.675 0.365 0.675 0.365 0.625 0.145 0.625 0.145 0.675 0.175 0.675 0.175 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01015 ;
  END A1N
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.635 0.635 0.495 0.665 0.495 0.665 0.425 0.415 0.425 0.415 0.475 0.58 0.475 0.58 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.045 0.835 0.905 0.905 0.905 0.905 0.325 0.7 0.325 0.7 0.185 0.65 0.185 0.65 0.375 0.85 0.375 0.85 0.855 0.785 0.855 0.785 1.045 ;
    END
    ANTENNADIFFAREA 0.07075 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 1 0.235 1 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.775 0.035 0.775 0.27 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.19 0.17 0.19 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.18 1.06 0.18 0.99 0.075 0.99 0.075 0.575 0.425 0.575 0.425 0.595 0.515 0.595 0.515 0.525 0.295 0.525 0.295 0.095 0.245 0.095 0.245 0.525 0.025 0.525 0.025 1.06 ;
      POLYGON 0.7 1.015 0.7 0.825 0.38 0.825 0.38 1.015 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1.015 ;
  END
END AOI2XB1_X1M_A12TUL_C35

MACRO NAND2XB_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2XB_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.565 0.175 0.565 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.008575 ;
  END BN
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.705 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0238 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.27 0.58 0.27 0.58 0.825 0.38 0.825 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.05775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.87 0.235 0.87 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.18 1.085 0.18 1.015 0.085 1.015 0.085 0.495 0.31 0.495 0.31 0.595 0.36 0.595 0.36 0.445 0.17 0.445 0.17 0.095 0.1 0.095 0.1 0.445 0.03 0.445 0.03 1.085 ;
  END
END NAND2XB_X1M_A12TUL_C35

MACRO OA1B2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA1B2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.235 0.725 0.235 0.525 0.165 0.525 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.805 0.505 0.805 0.505 0.525 0.435 0.525 0.435 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.105 0.71 1.005 0.77 1.005 0.77 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.715 0.375 0.715 0.925 0.64 0.925 0.64 1.105 ;
    END
    ANTENNADIFFAREA 0.07325 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.22 0.17 0.22 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.04 0.16 0.835 0.075 0.835 0.075 0.375 0.415 0.375 0.415 0.475 0.58 0.475 0.58 0.535 0.63 0.535 0.63 0.425 0.465 0.425 0.465 0.325 0.305 0.325 0.305 0.095 0.235 0.095 0.235 0.325 0.025 0.325 0.025 0.885 0.11 0.885 0.11 1.04 ;
  END
END OA1B2_X1M_A12TUL_C35

MACRO OR2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OR2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.565 0.17 0.565 0.17 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013825 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.305 0.475 0.305 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013825 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.045 0.565 0.905 0.635 0.905 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.045 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 0.17 0.18 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.05 0.16 0.86 0.075 0.86 0.075 0.375 0.445 0.375 0.445 0.57 0.495 0.57 0.495 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.325 0.025 0.325 0.025 0.91 0.11 0.91 0.11 1.05 ;
  END
END OR2_X0P7M_A12TUL_C35

MACRO AND2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.565 0.17 0.565 0.17 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0098 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0098 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.275 0.58 0.275 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.034875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0.17 1.165 0.17 1.025 0.1 1.025 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.305 1.105 0.305 0.875 0.495 0.875 0.495 0.325 0.16 0.325 0.16 0.13 0.11 0.13 0.11 0.375 0.445 0.375 0.445 0.825 0.255 0.825 0.255 1.015 0.235 1.015 0.235 1.105 ;
  END
END AND2_X0P5M_A12TUL_C35

MACRO OAI21B_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI21B_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.655 0.635 0.425 0.415 0.425 0.415 0.475 0.58 0.475 0.58 0.655 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.475 0.715 0.475 0.715 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.575 0.365 0.525 0.23 0.525 0.23 0.295 0.175 0.295 0.175 0.505 0.145 0.505 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00875 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.905 0.875 0.905 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.85 0.375 0.85 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.07675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.305 1.165 0.305 1.02 0.235 1.02 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.175 0.305 0.035 0.64 0.035 0.64 0.165 0.71 0.165 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.175 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.105 0.16 0.675 0.505 0.675 0.505 0.525 0.435 0.525 0.435 0.625 0.085 0.625 0.085 0.175 0.175 0.175 0.175 0.095 0.035 0.095 0.035 0.675 0.11 0.675 0.11 1.105 ;
      POLYGON 0.845 0.275 0.845 0.095 0.775 0.095 0.775 0.225 0.575 0.225 0.575 0.095 0.505 0.095 0.505 0.275 ;
  END
END OAI21B_X1M_A12TUL_C35

MACRO NAND4_X0P5A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND4_X0P5A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.495 0.435 0.495 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.595 0.31 0.595 0.31 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.175 0.475 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.115 0.575 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.235 0.925 0.235 1.115 0.305 1.115 0.305 0.975 0.505 0.975 0.505 1.115 ;
    END
    ANTENNADIFFAREA 0.03675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 1.04 0.37 1.04 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND4_X0P5A_A12TUL_C35

MACRO NOR4BB_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR4BB_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0084 ;
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.395 0.31 0.395 0.31 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0084 ;
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.775 0.64 0.565 0.57 0.565 0.57 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.635 0.505 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.435 0.495 0.435 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.105 0.845 1.005 0.905 1.005 0.905 0.225 0.85 0.225 0.85 0.085 0.77 0.085 0.77 0.225 0.575 0.225 0.575 0.09 0.505 0.09 0.505 0.275 0.85 0.275 0.85 0.925 0.775 0.925 0.775 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.185 0.44 0.035 0.64 0.035 0.64 0.165 0.71 0.165 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.185 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.31 1.105 0.31 1.025 0.28 1.025 0.28 0.875 0.765 0.875 0.765 0.665 0.715 0.665 0.715 0.825 0.085 0.825 0.085 0.175 0.19 0.175 0.19 0.125 0.035 0.125 0.035 0.875 0.23 0.875 0.23 1.105 ;
  END
END NOR4BB_X0P5M_A12TUL_C35

MACRO AND4_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND4_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.625 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.625 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.365 0.725 0.365 0.595 0.31 0.595 0.31 0.705 0.15 0.705 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.505 0.625 0.505 0.495 0.435 0.495 0.435 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.07 0.835 0.93 0.905 0.93 0.905 0.195 0.845 0.195 0.845 0.085 0.775 0.085 0.775 0.27 0.85 0.27 0.85 0.88 0.785 0.88 0.785 1.07 ;
    END
    ANTENNADIFFAREA 0.034875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.885 0.64 0.885 0.64 1.165 0.44 1.165 0.44 1.005 0.37 1.005 0.37 1.165 0.17 1.165 0.17 1.005 0.1 1.005 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.64 0.035 0.64 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.08 0.565 0.815 0.765 0.815 0.765 0.625 0.715 0.625 0.715 0.765 0.515 0.765 0.515 0.86 0.085 0.86 0.085 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.035 0.305 0.035 0.91 0.245 0.91 0.245 1.08 0.295 1.08 0.295 0.91 0.515 0.91 0.515 1.08 ;
  END
END AND4_X0P5M_A12TUL_C35

MACRO NAND4BB_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND4BB_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.725 0.235 0.575 0.365 0.575 0.365 0.525 0.145 0.525 0.145 0.575 0.165 0.575 0.165 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.665 0.31 0.665 0.31 0.805 0.15 0.805 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.675 0.645 0.425 0.415 0.425 0.415 0.475 0.565 0.475 0.565 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0175 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.565 0.435 0.565 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0175 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.11 0.845 0.975 0.905 0.975 0.905 0.195 0.845 0.195 0.845 0.09 0.775 0.09 0.775 0.27 0.85 0.27 0.85 0.925 0.505 0.925 0.505 1.105 0.575 1.105 0.575 0.975 0.775 0.975 0.775 1.11 ;
    END
    ANTENNADIFFAREA 0.0585 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 1.035 0.64 1.035 0.64 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.11 0.17 0.93 0.075 0.93 0.075 0.375 0.715 0.375 0.715 0.57 0.77 0.57 0.77 0.325 0.305 0.325 0.305 0.09 0.235 0.09 0.235 0.325 0.025 0.325 0.025 0.98 0.1 0.98 0.1 1.11 ;
  END
END NAND4BB_X0P7M_A12TUL_C35

MACRO BUFH_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUFH_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.525 0.145 0.525 0.145 0.575 0.345 0.575 0.345 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 0.84 0.565 0.84 0.605 0.91 0.605 0.91 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUFH_X4M_A12TL_C35

MACRO BUF_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUF_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0364 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.85 0.1 0.85 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.025 0.295 0.775 0.495 0.775 0.495 0.565 0.83 0.565 0.83 0.585 0.92 0.585 0.92 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.115 0.245 0.115 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 1.025 ;
  END
END BUF_X4M_A12TL_C35

MACRO INV_X3M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X3M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X3M_A12TH_C35

MACRO INV_X4B_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X4B_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.144 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.275 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.275 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X4B_A12TH_C35

MACRO INV_X5M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.161 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.85 0.375 0.85 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
END INV_X5M_A12TH_C35

MACRO INV_X0P8M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X0P8M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.058125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P8M_A12TH_C35

MACRO INV_X7P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X7P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.675 1.04 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.77 0.525 0.77 0.425 0.55 0.425 0.55 0.475 0.72 0.475 0.72 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2422 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.88 0.515 0.88 0.515 0.985 0.565 0.985 0.565 0.88 0.785 0.88 0.785 0.985 0.835 0.985 0.835 0.88 1.055 0.88 1.055 0.985 1.105 0.985 1.105 0.88 1.325 0.88 1.325 0.305 1.105 0.305 1.105 0.2 1.055 0.2 1.055 0.305 0.835 0.305 0.835 0.2 0.785 0.2 0.785 0.305 0.565 0.305 0.565 0.2 0.515 0.2 0.515 0.305 0.295 0.305 0.295 0.185 0.245 0.185 0.245 0.375 1.255 0.375 1.255 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.245 0.44 0.245 0.44 0.035 0.64 0.035 0.64 0.245 0.71 0.245 0.71 0.035 0.91 0.035 0.91 0.245 0.98 0.245 0.98 0.035 1.175 0.035 1.175 0.255 1.255 0.255 1.255 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
END INV_X7P5M_A12TH_C35

MACRO INV_X6M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X6M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.5 0.525 0.5 0.425 0.28 0.425 0.28 0.475 0.45 0.475 0.45 0.525 0.145 0.525 0.145 0.575 0.72 0.575 0.72 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1932 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.01 0.295 0.875 0.515 0.875 0.515 0.995 0.565 0.995 0.565 0.875 0.785 0.875 0.785 0.995 0.835 0.995 0.835 0.875 1.04 0.875 1.04 0.32 0.835 0.32 0.835 0.2 0.785 0.2 0.785 0.32 0.565 0.32 0.565 0.2 0.515 0.2 0.515 0.32 0.295 0.32 0.295 0.185 0.245 0.185 0.245 0.375 0.985 0.375 0.985 0.82 0.245 0.82 0.245 1.01 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
END INV_X6M_A12TH_C35

MACRO XOR3_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN XOR3_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 4.59 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 2.075 0.525 2.125 0.575 ;
        RECT 3.31 0.525 3.44 0.575 ;
      LAYER M1 ;
        RECT 2.06 0.43 2.14 0.645 ;
        POLYGON 3.48 0.655 3.48 0.525 3.27 0.525 3.27 0.655 3.34 0.655 3.34 0.575 3.41 0.575 3.41 0.655 ;
      LAYER M2 ;
        RECT 2.025 0.525 3.49 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 LAYER M1 ;
    ANTENNAGATEAREA 0.08995 LAYER M2 ;
    ANTENNAGATEAREA 0.08995 LAYER M3 ;
    ANTENNAGATEAREA 0.08995 LAYER M4 ;
    ANTENNAGATEAREA 0.08995 LAYER M5 ;
    ANTENNAGATEAREA 0.08995 LAYER M6 ;
    ANTENNAGATEAREA 0.08995 LAYER M7 ;
    ANTENNAGATEAREA 0.08995 LAYER M8 ;
    ANTENNAGATEAREA 0.08995 LAYER AP ;
    ANTENNAMAXAREACAR 0.5341615 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2018634 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.295 0.625 1.425 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 1.455 0.685 1.455 0.505 1.385 0.505 1.385 0.615 1.32 0.615 1.32 0.505 1.25 0.505 1.25 0.685 ;
        POLYGON 1.99 0.685 1.99 0.525 1.92 0.525 1.92 0.615 1.855 0.615 1.855 0.505 1.785 0.505 1.785 0.685 ;
      LAYER M2 ;
        RECT 1.245 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04165 LAYER M1 ;
    ANTENNAGATEAREA 0.09135 LAYER M2 ;
    ANTENNAGATEAREA 0.09135 LAYER M3 ;
    ANTENNAGATEAREA 0.09135 LAYER M4 ;
    ANTENNAGATEAREA 0.09135 LAYER M5 ;
    ANTENNAGATEAREA 0.09135 LAYER M6 ;
    ANTENNAGATEAREA 0.09135 LAYER M7 ;
    ANTENNAGATEAREA 0.09135 LAYER M8 ;
    ANTENNAGATEAREA 0.09135 LAYER AP ;
    ANTENNAMAXAREACAR 0.6806723 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1560625 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.675 0.665 0.625 0.465 0.625 0.465 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.067725 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 1.015 4.075 0.875 4.295 0.875 4.295 1.005 4.345 1.005 4.345 0.875 4.55 0.875 4.55 0.325 4.345 0.325 4.345 0.19 4.295 0.19 4.295 0.325 4.075 0.325 4.075 0.185 4.025 0.185 4.025 0.375 4.495 0.375 4.495 0.825 4.025 0.825 4.025 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
        RECT 3.485 1.175 3.535 1.225 ;
        RECT 3.62 1.175 3.67 1.225 ;
        RECT 3.755 1.175 3.805 1.225 ;
        RECT 3.89 1.175 3.94 1.225 ;
        RECT 4.025 1.175 4.075 1.225 ;
        RECT 4.16 1.175 4.21 1.225 ;
        RECT 4.295 1.175 4.345 1.225 ;
        RECT 4.43 1.175 4.48 1.225 ;
      LAYER M1 ;
        POLYGON 4.59 1.235 4.59 1.165 4.49 1.165 4.49 0.93 4.42 0.93 4.42 1.165 4.22 1.165 4.22 0.945 4.15 0.945 4.15 1.165 3.95 1.165 3.95 0.845 3.88 0.845 3.88 1.165 3.145 1.165 3.145 1.03 3.065 1.03 3.065 1.165 2.87 1.165 2.87 0.775 2.8 0.775 2.8 1.165 2.6 1.165 2.6 0.93 2.53 0.93 2.53 1.165 2.33 1.165 2.33 0.93 2.26 0.93 2.26 1.165 2.06 1.165 2.06 0.795 1.99 0.795 1.99 1.165 1.79 1.165 1.79 0.875 1.72 0.875 1.72 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 4.59 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
        RECT 3.485 -0.025 3.535 0.025 ;
        RECT 3.62 -0.025 3.67 0.025 ;
        RECT 3.755 -0.025 3.805 0.025 ;
        RECT 3.89 -0.025 3.94 0.025 ;
        RECT 4.025 -0.025 4.075 0.025 ;
        RECT 4.16 -0.025 4.21 0.025 ;
        RECT 4.295 -0.025 4.345 0.025 ;
        RECT 4.43 -0.025 4.48 0.025 ;
      LAYER M1 ;
        POLYGON 2.06 0.36 2.06 0.035 2.26 0.035 2.26 0.27 2.33 0.27 2.33 0.035 2.53 0.035 2.53 0.335 2.6 0.335 2.6 0.035 2.8 0.035 2.8 0.27 2.87 0.27 2.87 0.035 3.07 0.035 3.07 0.27 3.14 0.27 3.14 0.035 3.88 0.035 3.88 0.35 3.95 0.35 3.95 0.035 4.15 0.035 4.15 0.255 4.22 0.255 4.22 0.035 4.42 0.035 4.42 0.27 4.49 0.27 4.49 0.035 4.59 0.035 4.59 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.72 0.035 1.72 0.305 1.79 0.305 1.79 0.035 1.99 0.035 1.99 0.36 ;
      LAYER M2 ;
        RECT 0 -0.065 4.59 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.51 1.115 1.51 0.925 1.575 0.925 1.575 0.385 1.51 0.385 1.51 0.26 1.46 0.26 1.46 0.385 1.24 0.385 1.24 0.185 0.91 0.185 0.91 0.365 0.98 0.365 0.98 0.235 1.19 0.235 1.19 0.435 1.525 0.435 1.525 0.875 1.46 0.875 1.46 1.065 1.24 1.065 1.24 0.94 1.19 0.94 1.19 1.065 0.97 1.065 0.97 0.965 0.92 0.965 0.92 1.115 ;
      POLYGON 3.67 1.105 3.67 0.915 3.62 0.915 3.62 1.055 3.265 1.055 3.265 0.925 2.995 0.925 2.995 0.655 2.79 0.655 2.79 0.375 3.41 0.375 3.41 0.195 3.34 0.195 3.34 0.325 2.995 0.325 2.995 0.2 2.945 0.2 2.945 0.325 2.74 0.325 2.74 0.705 2.945 0.705 2.945 0.975 3.215 0.975 3.215 1.105 ;
      POLYGON 0.835 1.02 0.835 0.895 1.04 0.895 1.04 1.005 1.12 1.005 1.12 0.845 0.415 0.845 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.375 0.835 0.375 0.835 0.135 1.325 0.135 1.325 0.325 1.375 0.325 1.375 0.085 0.785 0.085 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.365 0.325 0.365 0.425 0.31 0.425 0.31 0.515 0.16 0.515 0.16 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.895 0.515 0.895 0.515 1.02 0.565 1.02 0.565 0.895 0.785 0.895 0.785 1.02 ;
      POLYGON 2.455 1.015 2.455 0.875 2.675 0.875 2.675 0.405 2.455 0.405 2.455 0.265 2.405 0.265 2.405 0.455 2.625 0.455 2.625 0.825 2.405 0.825 2.405 1.015 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 3.41 1.005 3.41 0.825 3.115 0.825 3.115 0.475 3.67 0.475 3.67 0.23 3.62 0.23 3.62 0.425 3.065 0.425 3.065 0.515 2.86 0.515 2.86 0.585 3.065 0.585 3.065 0.875 3.34 0.875 3.34 1.005 ;
      POLYGON 1.385 1.005 1.385 0.825 1.225 0.825 1.225 0.745 0.9 0.745 0.9 0.475 1.12 0.475 1.12 0.29 1.04 0.29 1.04 0.425 0.85 0.425 0.85 0.795 1.175 0.795 1.175 0.875 1.315 0.875 1.315 1.005 ;
      POLYGON 1.915 1 1.915 0.745 1.71 0.745 1.71 0.425 1.915 0.425 1.915 0.165 1.865 0.165 1.865 0.375 1.66 0.375 1.66 0.795 1.865 0.795 1.865 1 ;
      POLYGON 3.805 0.9 3.805 0.775 3.875 0.775 3.875 0.575 4.34 0.575 4.34 0.595 4.43 0.595 4.43 0.525 3.875 0.525 3.875 0.42 3.805 0.42 3.805 0.085 3.205 0.085 3.205 0.27 3.275 0.27 3.275 0.135 3.485 0.135 3.485 0.26 3.535 0.26 3.535 0.135 3.755 0.135 3.755 0.47 3.825 0.47 3.825 0.725 3.185 0.725 3.185 0.775 3.485 0.775 3.485 0.9 3.535 0.9 3.535 0.775 3.755 0.775 3.755 0.9 ;
      POLYGON 2.185 0.89 2.185 0.75 2.25 0.75 2.25 0.325 2.185 0.325 2.185 0.185 2.135 0.185 2.135 0.375 2.2 0.375 2.2 0.7 2.135 0.7 2.135 0.89 ;
      POLYGON 2.355 0.875 2.355 0.595 2.54 0.595 2.54 0.525 2.305 0.525 2.305 0.805 2.245 0.805 2.245 0.875 ;
      POLYGON 1.19 0.685 1.19 0.525 0.97 0.525 0.97 0.685 1.05 0.685 1.05 0.595 1.11 0.595 1.11 0.685 ;
      POLYGON 3.75 0.675 3.75 0.545 3.68 0.545 3.68 0.625 3.61 0.625 3.61 0.545 3.54 0.545 3.54 0.675 ;
    LAYER M2 ;
      RECT 2.455 0.825 3.285 0.875 ;
      RECT 1.475 0.825 2.375 0.875 ;
      RECT 0.075 0.825 1.395 0.875 ;
      RECT 2.15 0.625 3.76 0.675 ;
      RECT 0.965 0.525 1.76 0.575 ;
    LAYER VIA1 ;
      RECT 3.105 0.825 3.235 0.875 ;
      RECT 2.505 0.825 2.635 0.875 ;
      RECT 2.275 0.825 2.325 0.875 ;
      RECT 1.525 0.825 1.575 0.875 ;
      RECT 1.215 0.825 1.345 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 3.58 0.625 3.71 0.675 ;
      RECT 2.2 0.625 2.25 0.675 ;
      RECT 1.66 0.525 1.71 0.575 ;
      RECT 1.015 0.525 1.145 0.575 ;
  END
END XOR3_X4M_A12TL_C35

MACRO BUF_X6M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUF_X6M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05355 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.88 0.785 0.88 0.785 1 0.835 1 0.835 0.88 1.055 0.88 1.055 1 1.105 1 1.105 0.88 1.31 0.88 1.31 0.325 1.105 0.325 1.105 0.205 1.055 0.205 1.055 0.325 0.835 0.325 0.835 0.205 0.785 0.205 0.785 0.325 0.565 0.325 0.565 0.19 0.515 0.19 0.515 0.38 1.255 0.38 1.255 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.27 1.25 0.27 1.25 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 1.1 0.565 1.1 0.585 1.19 0.585 1.19 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUF_X6M_A12TL_C35

MACRO XNOR3_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 4.59 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 2.07 0.525 2.12 0.575 ;
        RECT 3.31 0.525 3.44 0.575 ;
      LAYER M1 ;
        RECT 2.055 0.43 2.135 0.645 ;
        POLYGON 3.48 0.655 3.48 0.525 3.27 0.525 3.27 0.655 3.34 0.655 3.34 0.575 3.41 0.575 3.41 0.655 ;
      LAYER M2 ;
        RECT 2.02 0.525 3.49 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 LAYER M1 ;
    ANTENNAGATEAREA 0.08995 LAYER M2 ;
    ANTENNAGATEAREA 0.08995 LAYER M3 ;
    ANTENNAGATEAREA 0.08995 LAYER M4 ;
    ANTENNAGATEAREA 0.08995 LAYER M5 ;
    ANTENNAGATEAREA 0.08995 LAYER M6 ;
    ANTENNAGATEAREA 0.08995 LAYER M7 ;
    ANTENNAGATEAREA 0.08995 LAYER M8 ;
    ANTENNAGATEAREA 0.08995 LAYER AP ;
    ANTENNAMAXAREACAR 0.5341615 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2018634 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.015 0.625 1.145 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 1.995 0.675 1.995 0.52 1.925 0.52 1.925 0.625 1.855 0.625 1.855 0.495 1.785 0.495 1.785 0.675 ;
        POLYGON 1.19 0.69 1.19 0.53 1.11 0.53 1.11 0.62 1.05 0.62 1.05 0.53 0.97 0.53 0.97 0.69 ;
      LAYER M2 ;
        RECT 0.965 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04165 LAYER M1 ;
    ANTENNAGATEAREA 0.09135 LAYER M2 ;
    ANTENNAGATEAREA 0.09135 LAYER M3 ;
    ANTENNAGATEAREA 0.09135 LAYER M4 ;
    ANTENNAGATEAREA 0.09135 LAYER M5 ;
    ANTENNAGATEAREA 0.09135 LAYER M6 ;
    ANTENNAGATEAREA 0.09135 LAYER M7 ;
    ANTENNAGATEAREA 0.09135 LAYER M8 ;
    ANTENNAGATEAREA 0.09135 LAYER AP ;
    ANTENNAMAXAREACAR 0.6470588 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1560625 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.465 0.625 0.465 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.067725 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 1.015 4.075 0.875 4.295 0.875 4.295 1.005 4.345 1.005 4.345 0.875 4.55 0.875 4.55 0.325 4.345 0.325 4.345 0.19 4.295 0.19 4.295 0.325 4.075 0.325 4.075 0.185 4.025 0.185 4.025 0.375 4.495 0.375 4.495 0.825 4.025 0.825 4.025 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
        RECT 3.485 1.175 3.535 1.225 ;
        RECT 3.62 1.175 3.67 1.225 ;
        RECT 3.755 1.175 3.805 1.225 ;
        RECT 3.89 1.175 3.94 1.225 ;
        RECT 4.025 1.175 4.075 1.225 ;
        RECT 4.16 1.175 4.21 1.225 ;
        RECT 4.295 1.175 4.345 1.225 ;
        RECT 4.43 1.175 4.48 1.225 ;
      LAYER M1 ;
        POLYGON 4.59 1.235 4.59 1.165 4.49 1.165 4.49 0.93 4.42 0.93 4.42 1.165 4.22 1.165 4.22 0.945 4.15 0.945 4.15 1.165 3.95 1.165 3.95 0.845 3.88 0.845 3.88 1.165 3.145 1.165 3.145 1.03 3.065 1.03 3.065 1.165 2.87 1.165 2.87 0.775 2.8 0.775 2.8 1.165 2.6 1.165 2.6 0.93 2.53 0.93 2.53 1.165 2.33 1.165 2.33 0.93 2.26 0.93 2.26 1.165 2.06 1.165 2.06 0.795 1.99 0.795 1.99 1.165 1.79 1.165 1.79 0.865 1.72 0.865 1.72 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 4.59 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
        RECT 3.485 -0.025 3.535 0.025 ;
        RECT 3.62 -0.025 3.67 0.025 ;
        RECT 3.755 -0.025 3.805 0.025 ;
        RECT 3.89 -0.025 3.94 0.025 ;
        RECT 4.025 -0.025 4.075 0.025 ;
        RECT 4.16 -0.025 4.21 0.025 ;
        RECT 4.295 -0.025 4.345 0.025 ;
        RECT 4.43 -0.025 4.48 0.025 ;
      LAYER M1 ;
        POLYGON 2.06 0.36 2.06 0.035 2.26 0.035 2.26 0.27 2.33 0.27 2.33 0.035 2.53 0.035 2.53 0.335 2.6 0.335 2.6 0.035 2.8 0.035 2.8 0.27 2.87 0.27 2.87 0.035 3.07 0.035 3.07 0.27 3.14 0.27 3.14 0.035 3.88 0.035 3.88 0.35 3.95 0.35 3.95 0.035 4.15 0.035 4.15 0.255 4.22 0.255 4.22 0.035 4.42 0.035 4.42 0.27 4.49 0.27 4.49 0.035 4.59 0.035 4.59 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.72 0.035 1.72 0.31 1.79 0.31 1.79 0.035 1.99 0.035 1.99 0.36 ;
      LAYER M2 ;
        RECT 0 -0.065 4.59 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.51 1.115 1.51 0.925 1.58 0.925 1.58 0.385 1.51 0.385 1.51 0.26 1.46 0.26 1.46 0.385 1.24 0.385 1.24 0.185 0.91 0.185 0.91 0.365 0.98 0.365 0.98 0.235 1.19 0.235 1.19 0.435 1.53 0.435 1.53 0.875 1.46 0.875 1.46 1.065 1.24 1.065 1.24 0.94 1.19 0.94 1.19 1.065 0.97 1.065 0.97 0.965 0.92 0.965 0.92 1.115 ;
      POLYGON 3.67 1.105 3.67 0.915 3.62 0.915 3.62 1.055 3.265 1.055 3.265 0.925 2.995 0.925 2.995 0.655 2.79 0.655 2.79 0.37 3.41 0.37 3.41 0.19 3.34 0.19 3.34 0.32 2.995 0.32 2.995 0.195 2.945 0.195 2.945 0.32 2.74 0.32 2.74 0.705 2.945 0.705 2.945 0.975 3.215 0.975 3.215 1.105 ;
      POLYGON 0.835 1.02 0.835 0.895 1.04 0.895 1.04 1.005 1.12 1.005 1.12 0.845 0.415 0.845 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.365 0.835 0.365 0.835 0.135 1.325 0.135 1.325 0.325 1.375 0.325 1.375 0.085 0.785 0.085 0.785 0.315 0.565 0.315 0.565 0.19 0.515 0.19 0.515 0.315 0.365 0.315 0.365 0.425 0.31 0.425 0.31 0.515 0.15 0.515 0.15 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.895 0.515 0.895 0.515 1.02 0.565 1.02 0.565 0.895 0.785 0.895 0.785 1.02 ;
      POLYGON 2.455 1.015 2.455 0.875 2.67 0.875 2.67 0.405 2.455 0.405 2.455 0.265 2.405 0.265 2.405 0.455 2.62 0.455 2.62 0.825 2.405 0.825 2.405 1.015 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 3.41 1.005 3.41 0.825 3.115 0.825 3.115 0.47 3.67 0.47 3.67 0.23 3.62 0.23 3.62 0.42 3.065 0.42 3.065 0.515 2.86 0.515 2.86 0.585 3.065 0.585 3.065 0.875 3.34 0.875 3.34 1.005 ;
      POLYGON 1.385 1.005 1.385 0.825 1.225 0.825 1.225 0.745 0.9 0.745 0.9 0.47 1.12 0.47 1.12 0.295 1.04 0.295 1.04 0.42 0.85 0.42 0.85 0.795 1.175 0.795 1.175 0.875 1.315 0.875 1.315 1.005 ;
      POLYGON 1.915 1 1.915 0.745 1.71 0.745 1.71 0.43 1.915 0.43 1.915 0.165 1.865 0.165 1.865 0.38 1.66 0.38 1.66 0.795 1.865 0.795 1.865 1 ;
      POLYGON 3.805 0.9 3.805 0.775 3.875 0.775 3.875 0.575 4.34 0.575 4.34 0.595 4.43 0.595 4.43 0.525 3.875 0.525 3.875 0.42 3.805 0.42 3.805 0.085 3.205 0.085 3.205 0.27 3.275 0.27 3.275 0.135 3.485 0.135 3.485 0.26 3.535 0.26 3.535 0.135 3.755 0.135 3.755 0.47 3.825 0.47 3.825 0.725 3.185 0.725 3.185 0.775 3.485 0.775 3.485 0.9 3.535 0.9 3.535 0.775 3.755 0.775 3.755 0.9 ;
      POLYGON 2.185 0.89 2.185 0.75 2.25 0.75 2.25 0.325 2.185 0.325 2.185 0.185 2.135 0.185 2.135 0.375 2.2 0.375 2.2 0.7 2.135 0.7 2.135 0.89 ;
      POLYGON 2.355 0.875 2.355 0.595 2.54 0.595 2.54 0.525 2.305 0.525 2.305 0.805 2.235 0.805 2.235 0.875 ;
      POLYGON 1.455 0.695 1.455 0.515 1.25 0.515 1.25 0.695 1.32 0.695 1.32 0.585 1.385 0.585 1.385 0.695 ;
      POLYGON 3.75 0.675 3.75 0.545 3.68 0.545 3.68 0.625 3.61 0.625 3.61 0.545 3.54 0.545 3.54 0.675 ;
    LAYER M2 ;
      RECT 2.45 0.825 3.295 0.875 ;
      RECT 1.48 0.825 2.37 0.875 ;
      RECT 0.075 0.825 1.395 0.875 ;
      RECT 2.15 0.625 3.76 0.675 ;
      RECT 1.235 0.525 1.76 0.575 ;
    LAYER VIA1 ;
      RECT 3.115 0.825 3.245 0.875 ;
      RECT 2.5 0.825 2.63 0.875 ;
      RECT 2.27 0.825 2.32 0.875 ;
      RECT 1.53 0.825 1.58 0.875 ;
      RECT 1.215 0.825 1.345 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 3.58 0.625 3.71 0.675 ;
      RECT 2.2 0.625 2.25 0.675 ;
      RECT 1.66 0.525 1.71 0.575 ;
      RECT 1.285 0.525 1.415 0.575 ;
  END
END XNOR3_X4M_A12TL_C35

MACRO INV_X4M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X4M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X4M_A12TH_C35

MACRO XNOR3_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 4.59 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 2.07 0.525 2.12 0.575 ;
        RECT 3.31 0.525 3.44 0.575 ;
      LAYER M1 ;
        RECT 2.055 0.43 2.135 0.645 ;
        POLYGON 3.48 0.655 3.48 0.525 3.27 0.525 3.27 0.655 3.34 0.655 3.34 0.575 3.41 0.575 3.41 0.655 ;
      LAYER M2 ;
        RECT 2.02 0.525 3.49 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 LAYER M1 ;
    ANTENNAGATEAREA 0.08995 LAYER M2 ;
    ANTENNAGATEAREA 0.08995 LAYER M3 ;
    ANTENNAGATEAREA 0.08995 LAYER M4 ;
    ANTENNAGATEAREA 0.08995 LAYER M5 ;
    ANTENNAGATEAREA 0.08995 LAYER M6 ;
    ANTENNAGATEAREA 0.08995 LAYER M7 ;
    ANTENNAGATEAREA 0.08995 LAYER M8 ;
    ANTENNAGATEAREA 0.08995 LAYER AP ;
    ANTENNAMAXAREACAR 0.5341615 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2018634 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.015 0.625 1.145 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 1.995 0.675 1.995 0.52 1.925 0.52 1.925 0.625 1.855 0.625 1.855 0.495 1.785 0.495 1.785 0.675 ;
        POLYGON 1.19 0.69 1.19 0.53 1.11 0.53 1.11 0.62 1.05 0.62 1.05 0.53 0.97 0.53 0.97 0.69 ;
      LAYER M2 ;
        RECT 0.965 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04165 LAYER M1 ;
    ANTENNAGATEAREA 0.09135 LAYER M2 ;
    ANTENNAGATEAREA 0.09135 LAYER M3 ;
    ANTENNAGATEAREA 0.09135 LAYER M4 ;
    ANTENNAGATEAREA 0.09135 LAYER M5 ;
    ANTENNAGATEAREA 0.09135 LAYER M6 ;
    ANTENNAGATEAREA 0.09135 LAYER M7 ;
    ANTENNAGATEAREA 0.09135 LAYER M8 ;
    ANTENNAGATEAREA 0.09135 LAYER AP ;
    ANTENNAMAXAREACAR 0.6470588 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1560625 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.465 0.625 0.465 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.067725 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 1.015 4.075 0.875 4.295 0.875 4.295 1.005 4.345 1.005 4.345 0.875 4.55 0.875 4.55 0.325 4.345 0.325 4.345 0.19 4.295 0.19 4.295 0.325 4.075 0.325 4.075 0.185 4.025 0.185 4.025 0.375 4.495 0.375 4.495 0.825 4.025 0.825 4.025 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
        RECT 3.485 1.175 3.535 1.225 ;
        RECT 3.62 1.175 3.67 1.225 ;
        RECT 3.755 1.175 3.805 1.225 ;
        RECT 3.89 1.175 3.94 1.225 ;
        RECT 4.025 1.175 4.075 1.225 ;
        RECT 4.16 1.175 4.21 1.225 ;
        RECT 4.295 1.175 4.345 1.225 ;
        RECT 4.43 1.175 4.48 1.225 ;
      LAYER M1 ;
        POLYGON 4.59 1.235 4.59 1.165 4.49 1.165 4.49 0.93 4.42 0.93 4.42 1.165 4.22 1.165 4.22 0.945 4.15 0.945 4.15 1.165 3.95 1.165 3.95 0.845 3.88 0.845 3.88 1.165 3.145 1.165 3.145 1.03 3.065 1.03 3.065 1.165 2.87 1.165 2.87 0.775 2.8 0.775 2.8 1.165 2.6 1.165 2.6 0.93 2.53 0.93 2.53 1.165 2.33 1.165 2.33 0.93 2.26 0.93 2.26 1.165 2.06 1.165 2.06 0.795 1.99 0.795 1.99 1.165 1.79 1.165 1.79 0.865 1.72 0.865 1.72 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 4.59 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
        RECT 3.485 -0.025 3.535 0.025 ;
        RECT 3.62 -0.025 3.67 0.025 ;
        RECT 3.755 -0.025 3.805 0.025 ;
        RECT 3.89 -0.025 3.94 0.025 ;
        RECT 4.025 -0.025 4.075 0.025 ;
        RECT 4.16 -0.025 4.21 0.025 ;
        RECT 4.295 -0.025 4.345 0.025 ;
        RECT 4.43 -0.025 4.48 0.025 ;
      LAYER M1 ;
        POLYGON 2.06 0.36 2.06 0.035 2.26 0.035 2.26 0.27 2.33 0.27 2.33 0.035 2.53 0.035 2.53 0.335 2.6 0.335 2.6 0.035 2.8 0.035 2.8 0.27 2.87 0.27 2.87 0.035 3.07 0.035 3.07 0.27 3.14 0.27 3.14 0.035 3.88 0.035 3.88 0.35 3.95 0.35 3.95 0.035 4.15 0.035 4.15 0.255 4.22 0.255 4.22 0.035 4.42 0.035 4.42 0.27 4.49 0.27 4.49 0.035 4.59 0.035 4.59 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.72 0.035 1.72 0.31 1.79 0.31 1.79 0.035 1.99 0.035 1.99 0.36 ;
      LAYER M2 ;
        RECT 0 -0.065 4.59 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.51 1.115 1.51 0.925 1.58 0.925 1.58 0.385 1.51 0.385 1.51 0.26 1.46 0.26 1.46 0.385 1.24 0.385 1.24 0.185 0.91 0.185 0.91 0.365 0.98 0.365 0.98 0.235 1.19 0.235 1.19 0.435 1.53 0.435 1.53 0.875 1.46 0.875 1.46 1.065 1.24 1.065 1.24 0.94 1.19 0.94 1.19 1.065 0.97 1.065 0.97 0.965 0.92 0.965 0.92 1.115 ;
      POLYGON 3.67 1.105 3.67 0.915 3.62 0.915 3.62 1.055 3.265 1.055 3.265 0.925 2.995 0.925 2.995 0.655 2.79 0.655 2.79 0.37 3.41 0.37 3.41 0.19 3.34 0.19 3.34 0.32 2.995 0.32 2.995 0.195 2.945 0.195 2.945 0.32 2.74 0.32 2.74 0.705 2.945 0.705 2.945 0.975 3.215 0.975 3.215 1.105 ;
      POLYGON 0.835 1.02 0.835 0.895 1.04 0.895 1.04 1.005 1.12 1.005 1.12 0.845 0.415 0.845 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.365 0.835 0.365 0.835 0.135 1.325 0.135 1.325 0.325 1.375 0.325 1.375 0.085 0.785 0.085 0.785 0.315 0.565 0.315 0.565 0.19 0.515 0.19 0.515 0.315 0.365 0.315 0.365 0.425 0.31 0.425 0.31 0.515 0.15 0.515 0.15 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.895 0.515 0.895 0.515 1.02 0.565 1.02 0.565 0.895 0.785 0.895 0.785 1.02 ;
      POLYGON 2.455 1.015 2.455 0.875 2.67 0.875 2.67 0.405 2.455 0.405 2.455 0.265 2.405 0.265 2.405 0.455 2.62 0.455 2.62 0.825 2.405 0.825 2.405 1.015 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 3.41 1.005 3.41 0.825 3.115 0.825 3.115 0.47 3.67 0.47 3.67 0.23 3.62 0.23 3.62 0.42 3.065 0.42 3.065 0.515 2.86 0.515 2.86 0.585 3.065 0.585 3.065 0.875 3.34 0.875 3.34 1.005 ;
      POLYGON 1.385 1.005 1.385 0.825 1.225 0.825 1.225 0.745 0.9 0.745 0.9 0.47 1.12 0.47 1.12 0.295 1.04 0.295 1.04 0.42 0.85 0.42 0.85 0.795 1.175 0.795 1.175 0.875 1.315 0.875 1.315 1.005 ;
      POLYGON 1.915 1 1.915 0.745 1.71 0.745 1.71 0.43 1.915 0.43 1.915 0.165 1.865 0.165 1.865 0.38 1.66 0.38 1.66 0.795 1.865 0.795 1.865 1 ;
      POLYGON 3.805 0.9 3.805 0.775 3.875 0.775 3.875 0.575 4.34 0.575 4.34 0.595 4.43 0.595 4.43 0.525 3.875 0.525 3.875 0.42 3.805 0.42 3.805 0.085 3.205 0.085 3.205 0.27 3.275 0.27 3.275 0.135 3.485 0.135 3.485 0.26 3.535 0.26 3.535 0.135 3.755 0.135 3.755 0.47 3.825 0.47 3.825 0.725 3.185 0.725 3.185 0.775 3.485 0.775 3.485 0.9 3.535 0.9 3.535 0.775 3.755 0.775 3.755 0.9 ;
      POLYGON 2.185 0.89 2.185 0.75 2.25 0.75 2.25 0.325 2.185 0.325 2.185 0.185 2.135 0.185 2.135 0.375 2.2 0.375 2.2 0.7 2.135 0.7 2.135 0.89 ;
      POLYGON 2.355 0.875 2.355 0.595 2.54 0.595 2.54 0.525 2.305 0.525 2.305 0.805 2.235 0.805 2.235 0.875 ;
      POLYGON 1.455 0.695 1.455 0.515 1.25 0.515 1.25 0.695 1.32 0.695 1.32 0.585 1.385 0.585 1.385 0.695 ;
      POLYGON 3.75 0.675 3.75 0.545 3.68 0.545 3.68 0.625 3.61 0.625 3.61 0.545 3.54 0.545 3.54 0.675 ;
    LAYER M2 ;
      RECT 2.45 0.825 3.295 0.875 ;
      RECT 1.48 0.825 2.37 0.875 ;
      RECT 0.075 0.825 1.395 0.875 ;
      RECT 2.15 0.625 3.76 0.675 ;
      RECT 1.235 0.525 1.76 0.575 ;
    LAYER VIA1 ;
      RECT 3.115 0.825 3.245 0.875 ;
      RECT 2.5 0.825 2.63 0.875 ;
      RECT 2.27 0.825 2.32 0.875 ;
      RECT 1.53 0.825 1.58 0.875 ;
      RECT 1.215 0.825 1.345 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 3.58 0.625 3.71 0.675 ;
      RECT 2.2 0.625 2.25 0.675 ;
      RECT 1.66 0.525 1.71 0.575 ;
      RECT 1.285 0.525 1.415 0.575 ;
  END
END XNOR3_X4M_A12TUL_C35

MACRO INV_X11M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X11M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.755 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.58 0.675 1.58 0.495 1.53 0.495 1.53 0.525 1.175 0.525 1.175 0.425 0.955 0.425 0.955 0.475 1.125 0.475 1.125 0.525 0.635 0.525 0.635 0.425 0.415 0.425 0.415 0.475 0.585 0.475 0.585 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 0.365 0.675 0.365 0.575 0.855 0.575 0.855 0.625 0.685 0.625 0.685 0.675 0.905 0.675 0.905 0.575 1.53 0.575 1.53 0.625 1.36 0.625 1.36 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3542 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.905 0.515 0.905 0.515 0.985 0.565 0.985 0.565 0.905 0.785 0.905 0.785 0.985 0.835 0.985 0.835 0.905 1.055 0.905 1.055 0.985 1.105 0.985 1.105 0.905 1.325 0.905 1.325 0.985 1.375 0.985 1.375 0.905 1.595 0.905 1.595 0.985 1.645 0.985 1.645 0.905 1.73 0.905 1.73 0.28 1.645 0.28 1.645 0.2 1.595 0.2 1.595 0.28 1.375 0.28 1.375 0.2 1.325 0.2 1.325 0.28 1.105 0.28 1.105 0.2 1.055 0.2 1.055 0.28 0.835 0.28 0.835 0.2 0.785 0.2 0.785 0.28 0.565 0.28 0.565 0.2 0.515 0.2 0.515 0.28 0.295 0.28 0.295 0.185 0.245 0.185 0.245 0.375 1.635 0.375 1.635 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
      LAYER M1 ;
        POLYGON 1.755 1.235 1.755 1.165 1.525 1.165 1.525 0.955 1.445 0.955 1.445 1.165 1.255 1.165 1.255 0.955 1.175 0.955 1.175 1.165 0.985 1.165 0.985 0.955 0.905 0.955 0.905 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.755 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.365 0.035 0.365 0.23 0.445 0.23 0.445 0.035 0.635 0.035 0.635 0.23 0.715 0.23 0.715 0.035 0.905 0.035 0.905 0.23 0.985 0.23 0.985 0.035 1.175 0.035 1.175 0.23 1.255 0.23 1.255 0.035 1.445 0.035 1.445 0.23 1.525 0.23 1.525 0.035 1.755 0.035 1.755 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.755 0.065 ;
    END
  END VSS
END INV_X11M_A12TH_C35

MACRO BUFH_X2M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUFH_X2M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.595 0.515 0.595 0.515 0.525 0.425 0.525 0.425 0.535 0.28 0.535 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X2M_A12TL_C35

MACRO INV_X9M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X9M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.575 1.255 0.575 1.255 0.605 1.31 0.605 1.31 0.495 1.255 0.495 1.255 0.525 0.905 0.525 0.905 0.425 0.685 0.425 0.685 0.475 0.855 0.475 0.855 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 0.635 0.675 0.635 0.575 1.125 0.575 1.125 0.625 0.955 0.625 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2898 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.89 0.515 0.89 0.515 0.985 0.565 0.985 0.565 0.89 0.785 0.89 0.785 0.985 0.835 0.985 0.835 0.89 1.055 0.89 1.055 0.985 1.105 0.985 1.105 0.89 1.325 0.89 1.325 0.985 1.375 0.985 1.375 0.89 1.46 0.89 1.46 0.295 1.375 0.295 1.375 0.195 1.325 0.195 1.325 0.295 1.105 0.295 1.105 0.2 1.055 0.2 1.055 0.295 0.835 0.295 0.835 0.2 0.785 0.2 0.785 0.295 0.565 0.295 0.565 0.2 0.515 0.2 0.515 0.295 0.295 0.295 0.295 0.185 0.245 0.185 0.245 0.375 1.38 0.375 1.38 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.437 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 1.255 1.165 1.255 0.955 1.175 0.955 1.175 1.165 0.985 1.165 0.985 0.955 0.905 0.955 0.905 1.165 0.715 1.165 0.715 0.955 0.635 0.955 0.635 1.165 0.445 1.165 0.445 0.955 0.365 0.955 0.365 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.365 0.035 0.365 0.235 0.445 0.235 0.445 0.035 0.635 0.035 0.635 0.235 0.715 0.235 0.715 0.035 0.905 0.035 0.905 0.235 0.985 0.235 0.985 0.035 1.175 0.035 1.175 0.235 1.255 0.235 1.255 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
END INV_X9M_A12TH_C35

MACRO BUF_X9M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUF_X9M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.08085 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.99 0.7 0.88 0.92 0.88 0.92 0.975 0.97 0.975 0.97 0.88 1.19 0.88 1.19 0.975 1.24 0.975 1.24 0.88 1.46 0.88 1.46 0.975 1.51 0.975 1.51 0.88 1.73 0.88 1.73 0.975 1.78 0.975 1.78 0.88 1.865 0.88 1.865 0.32 1.78 0.32 1.78 0.22 1.73 0.22 1.73 0.32 1.51 0.32 1.51 0.225 1.46 0.225 1.46 0.32 1.24 0.32 1.24 0.225 1.19 0.225 1.19 0.32 0.97 0.32 0.97 0.225 0.92 0.225 0.92 0.32 0.7 0.32 0.7 0.21 0.65 0.21 0.65 0.4 1.785 0.4 1.785 0.8 0.65 0.8 0.65 0.99 ;
    END
    ANTENNADIFFAREA 0.437 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.655 1.165 1.655 0.945 1.585 0.945 1.585 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.945 1.045 0.945 1.045 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.355 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.585 0.035 1.585 0.255 1.655 0.255 1.655 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1 0.43 0.875 0.565 0.875 0.565 0.725 0.63 0.725 0.63 0.565 1.65 0.565 1.65 0.605 1.72 0.605 1.72 0.515 0.58 0.515 0.58 0.675 0.515 0.675 0.515 0.825 0.085 0.825 0.085 0.375 0.43 0.375 0.43 0.185 0.38 0.185 0.38 0.325 0.16 0.325 0.16 0.2 0.11 0.2 0.11 0.325 0.035 0.325 0.035 0.875 0.11 0.875 0.11 1 0.16 1 0.16 0.875 0.38 0.875 0.38 1 ;
  END
END BUF_X9M_A12TL_C35

MACRO INV_X1P2M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X1P2M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0385 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.13 0.245 0.13 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.055 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.305 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P2M_A12TH_C35

MACRO INV_X1P4M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X1P4M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.175 0.245 0.175 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P4M_A12TH_C35

MACRO XNOR3_X3M_A12TL_C35
  CLASS CORE ;
  FOREIGN XNOR3_X3M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.51 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.795 0.625 1.845 0.675 ;
        RECT 2.785 0.625 2.835 0.675 ;
      LAYER M1 ;
        POLYGON 2.91 0.675 2.91 0.605 2.815 0.605 2.815 0.515 2.735 0.515 2.735 0.675 ;
        RECT 1.785 0.42 1.855 0.71 ;
      LAYER M2 ;
        RECT 1.745 0.625 2.885 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 LAYER M1 ;
    ANTENNAGATEAREA 0.05495 LAYER M2 ;
    ANTENNAGATEAREA 0.05495 LAYER M3 ;
    ANTENNAGATEAREA 0.05495 LAYER M4 ;
    ANTENNAGATEAREA 0.05495 LAYER M5 ;
    ANTENNAGATEAREA 0.05495 LAYER M6 ;
    ANTENNAGATEAREA 0.05495 LAYER M7 ;
    ANTENNAGATEAREA 0.05495 LAYER M8 ;
    ANTENNAGATEAREA 0.05495 LAYER AP ;
    ANTENNAMAXAREACAR 0.8923078 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1098901 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.88 0.525 1.01 0.575 ;
        RECT 1.66 0.525 1.71 0.575 ;
      LAYER M1 ;
        POLYGON 1.05 0.65 1.05 0.525 0.84 0.525 0.84 0.65 0.91 0.65 0.91 0.575 0.98 0.575 0.98 0.65 ;
        RECT 1.65 0.42 1.72 0.71 ;
      LAYER M2 ;
        RECT 0.83 0.525 1.76 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0308 LAYER M1 ;
    ANTENNAGATEAREA 0.0924 LAYER M2 ;
    ANTENNAGATEAREA 0.0924 LAYER M3 ;
    ANTENNAGATEAREA 0.0924 LAYER M4 ;
    ANTENNAGATEAREA 0.0924 LAYER M5 ;
    ANTENNAGATEAREA 0.0924 LAYER M6 ;
    ANTENNAGATEAREA 0.0924 LAYER M7 ;
    ANTENNAGATEAREA 0.0924 LAYER M8 ;
    ANTENNAGATEAREA 0.0924 LAYER AP ;
    ANTENNAMAXAREACAR 0.659091 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.211039 LAYER VIA1 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.465 0.625 0.465 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.415 0.525 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05775 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 3.13 1.015 3.13 0.875 3.35 0.875 3.35 1 3.4 1 3.4 0.875 3.47 0.875 3.47 0.325 3.4 0.325 3.4 0.2 3.35 0.2 3.35 0.325 3.13 0.325 3.13 0.185 3.08 0.185 3.08 0.375 3.415 0.375 3.415 0.825 3.08 0.825 3.08 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
        RECT 3.35 1.175 3.4 1.225 ;
      LAYER M1 ;
        POLYGON 3.51 1.235 3.51 1.165 3.275 1.165 3.275 0.945 3.205 0.945 3.205 1.165 3.005 1.165 3.005 0.845 2.935 0.845 2.935 1.165 2.47 1.165 2.47 1.03 2.39 1.03 2.39 1.165 2.195 1.165 2.195 0.905 2.125 0.905 2.125 1.165 1.79 1.165 1.79 0.78 1.72 0.78 1.72 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.925 0.1 0.925 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.51 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
        RECT 3.35 -0.025 3.4 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.35 1.79 0.035 2.12 0.035 2.12 0.26 2.2 0.26 2.2 0.035 2.39 0.035 2.39 0.26 2.47 0.26 2.47 0.035 2.93 0.035 2.93 0.26 3.01 0.26 3.01 0.035 3.205 0.035 3.205 0.255 3.275 0.255 3.275 0.035 3.51 0.035 3.51 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.635 0.035 0.635 0.26 0.715 0.26 0.715 0.035 1.72 0.035 1.72 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 3.51 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.375 1.115 1.375 0.925 1.445 0.925 1.445 0.325 1.375 0.325 1.375 0.09 0.785 0.09 0.785 0.24 0.835 0.24 0.835 0.14 1.04 0.14 1.04 0.26 1.12 0.26 1.12 0.14 1.325 0.14 1.325 0.375 1.395 0.375 1.395 0.875 1.325 0.875 1.325 1.065 1.105 1.065 1.105 0.94 1.055 0.94 1.055 1.065 0.845 1.065 0.845 0.93 0.775 0.93 0.775 1.115 ;
      POLYGON 2.86 1.035 2.86 0.845 2.81 0.845 2.81 0.985 2.59 0.985 2.59 0.925 2.32 0.925 2.32 0.785 2.115 0.785 2.115 0.36 2.59 0.36 2.59 0.17 2.54 0.17 2.54 0.31 2.32 0.31 2.32 0.185 2.27 0.185 2.27 0.31 2.065 0.31 2.065 0.835 2.27 0.835 2.27 0.975 2.54 0.975 2.54 1.035 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
      POLYGON 1.25 1.005 1.25 0.825 1.09 0.825 1.09 0.725 0.775 0.725 0.775 0.465 1 0.465 1 0.415 0.725 0.415 0.725 0.775 1.04 0.775 1.04 0.875 1.18 0.875 1.18 1.005 ;
      POLYGON 0.98 1.005 0.98 0.825 0.415 0.825 0.415 0.725 0.36 0.725 0.36 0.475 0.415 0.475 0.415 0.36 1.255 0.36 1.255 0.2 1.175 0.2 1.175 0.31 0.565 0.31 0.565 0.185 0.515 0.185 0.515 0.31 0.365 0.31 0.365 0.425 0.31 0.425 0.31 0.515 0.16 0.515 0.16 0.585 0.31 0.585 0.31 0.775 0.365 0.775 0.365 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.91 0.875 0.91 1.005 ;
      POLYGON 1.915 0.995 1.915 0.855 1.98 0.855 1.98 0.3 1.915 0.3 1.915 0.16 1.865 0.16 1.865 0.35 1.93 0.35 1.93 0.805 1.865 0.805 1.865 0.995 ;
      POLYGON 1.645 0.97 1.645 0.78 1.575 0.78 1.575 0.35 1.645 0.35 1.645 0.16 1.595 0.16 1.595 0.3 1.525 0.3 1.525 0.83 1.595 0.83 1.595 0.97 ;
      POLYGON 2.725 0.915 2.725 0.775 3.02 0.775 3.02 0.585 3.35 0.585 3.35 0.515 3.02 0.515 3.02 0.31 2.725 0.31 2.725 0.17 2.675 0.17 2.675 0.36 2.97 0.36 2.97 0.725 2.675 0.725 2.675 0.915 ;
      POLYGON 2.6 0.875 2.6 0.665 2.385 0.665 2.385 0.46 2.89 0.46 2.89 0.41 2.335 0.41 2.335 0.515 2.185 0.515 2.185 0.585 2.335 0.585 2.335 0.715 2.54 0.715 2.54 0.825 2.39 0.825 2.39 0.875 ;
      POLYGON 1.32 0.675 1.32 0.52 1.25 0.52 1.25 0.625 1.18 0.625 1.18 0.52 1.11 0.52 1.11 0.675 ;
      RECT 2.44 0.52 2.675 0.6 ;
    LAYER M2 ;
      RECT 1.345 0.825 2.61 0.875 ;
      RECT 0.075 0.825 1.26 0.875 ;
      RECT 1.1 0.625 1.625 0.675 ;
      RECT 1.88 0.525 2.66 0.575 ;
    LAYER VIA1 ;
      RECT 2.43 0.825 2.56 0.875 ;
      RECT 1.395 0.825 1.445 0.875 ;
      RECT 1.08 0.825 1.21 0.875 ;
      RECT 0.125 0.825 0.255 0.875 ;
      RECT 1.525 0.625 1.575 0.675 ;
      RECT 1.15 0.625 1.28 0.675 ;
      RECT 2.48 0.525 2.61 0.575 ;
      RECT 1.93 0.525 1.98 0.575 ;
  END
END XNOR3_X3M_A12TL_C35

MACRO INV_X16M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X16M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.12 0.675 2.12 0.58 2.18 0.58 2.18 0.6 2.27 0.6 2.27 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 1.04 0.675 1.04 0.575 1.53 0.575 1.53 0.625 1.36 0.625 1.36 0.675 1.58 0.675 1.58 0.575 2.07 0.575 2.07 0.625 1.9 0.625 1.9 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5152 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 0.935 0.295 0.885 0.515 0.885 0.515 0.93 0.565 0.93 0.565 0.885 0.785 0.885 0.785 0.93 0.835 0.93 0.835 0.885 1.055 0.885 1.055 0.93 1.105 0.93 1.105 0.885 1.325 0.885 1.325 0.93 1.375 0.93 1.375 0.885 1.595 0.885 1.595 0.93 1.645 0.93 1.645 0.885 1.865 0.885 1.865 0.93 1.915 0.93 1.915 0.885 2.135 0.885 2.135 0.93 2.185 0.93 2.185 0.885 2.46 0.885 2.46 0.315 2.185 0.315 2.185 0.27 2.135 0.27 2.135 0.315 1.915 0.315 1.915 0.27 1.865 0.27 1.865 0.315 1.645 0.315 1.645 0.27 1.595 0.27 1.595 0.315 1.375 0.315 1.375 0.27 1.325 0.27 1.325 0.315 1.105 0.315 1.105 0.27 1.055 0.27 1.055 0.315 0.835 0.315 0.835 0.27 0.785 0.27 0.785 0.315 0.565 0.315 0.565 0.27 0.515 0.27 0.515 0.315 0.295 0.315 0.295 0.265 0.245 0.265 0.245 0.455 2.325 0.455 2.325 0.745 0.245 0.745 0.245 0.935 ;
    END
    ANTENNADIFFAREA 0.736 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
      LAYER M1 ;
        POLYGON 2.565 1.235 2.565 1.165 2.465 1.165 2.465 0.995 2.395 0.995 2.395 1.165 2.33 1.165 2.33 0.945 2.26 0.945 2.26 1.165 2.06 1.165 2.06 0.945 1.99 0.945 1.99 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.565 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 1.72 0.035 1.72 0.255 1.79 0.255 1.79 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.26 0.035 2.26 0.255 2.33 0.255 2.33 0.035 2.395 0.035 2.395 0.205 2.465 0.205 2.465 0.035 2.565 0.035 2.565 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 2.565 0.065 ;
    END
  END VSS
END INV_X16M_A12TL_C35

MACRO INV_X1P7M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X1P7M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05425 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.0775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P7M_A12TH_C35

MACRO INV_X2M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X2M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X2M_A12TH_C35

MACRO INV_X0P6M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X0P6M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01925 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.065 0.295 0.925 0.365 0.925 0.365 0.26 0.295 0.26 0.295 0.12 0.245 0.12 0.245 0.31 0.31 0.31 0.31 0.875 0.245 0.875 0.245 1.065 ;
    END
    ANTENNADIFFAREA 0.04125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.875 0.1 0.875 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.3 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.3 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P6M_A12TH_C35

MACRO INV_X1P2B_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X1P2B_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.225 0.295 0.225 0.295 0.095 0.245 0.095 0.245 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.043 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.18 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P2B_A12TH_C35

MACRO INV_X0P7M_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X0P7M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P7M_A12TH_C35

MACRO XOR2_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN XOR2_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.7 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.94 0.625 2.07 0.675 ;
        RECT 2.36 0.625 2.49 0.675 ;
      LAYER M1 ;
        POLYGON 2.12 0.675 2.12 0.565 2.07 0.565 2.07 0.625 1.985 0.625 1.985 0.565 1.935 0.565 1.935 0.625 1.85 0.625 1.85 0.565 1.8 0.565 1.8 0.675 ;
        POLYGON 2.52 0.685 2.52 0.495 2.47 0.495 2.47 0.615 2.385 0.615 2.385 0.495 2.33 0.495 2.33 0.685 ;
      LAYER M2 ;
        RECT 1.89 0.625 2.54 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 LAYER M1 ;
    ANTENNAGATEAREA 0.13545 LAYER M2 ;
    ANTENNAGATEAREA 0.13545 LAYER M3 ;
    ANTENNAGATEAREA 0.13545 LAYER M4 ;
    ANTENNAGATEAREA 0.13545 LAYER M5 ;
    ANTENNAGATEAREA 0.13545 LAYER M6 ;
    ANTENNAGATEAREA 0.13545 LAYER M7 ;
    ANTENNAGATEAREA 0.13545 LAYER M8 ;
    ANTENNAGATEAREA 0.13545 LAYER AP ;
    ANTENNAMAXAREACAR 0.560606 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1406928 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 1.205 0.575 1.205 0.425 0.985 0.425 0.985 0.475 1.155 0.475 1.155 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.05 1 2.05 0.875 2.255 0.875 2.255 0.325 2.05 0.325 2.05 0.2 2 0.2 2 0.325 1.78 0.325 1.78 0.185 1.45 0.185 1.45 0.365 1.52 0.365 1.52 0.235 1.73 0.235 1.73 0.375 2.2 0.375 2.2 0.825 1.915 0.825 1.915 0.725 1.43 0.725 1.43 0.775 1.865 0.775 1.865 0.875 2 0.875 2 1 ;
    END
    ANTENNADIFFAREA 0.255 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
      LAYER M1 ;
        POLYGON 2.7 1.235 2.7 1.165 2.6 1.165 2.6 0.875 2.53 0.875 2.53 1.165 2.33 1.165 2.33 0.925 2.26 0.925 2.26 1.165 1.255 1.165 1.255 1.03 1.175 1.03 1.175 1.165 0.98 1.165 0.98 0.845 0.91 0.845 0.91 1.165 0.71 1.165 0.71 0.845 0.64 0.845 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.7 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.18 1.25 0.18 1.25 0.035 2.26 0.035 2.26 0.275 2.33 0.275 2.33 0.035 2.53 0.035 2.53 0.305 2.6 0.305 2.6 0.035 2.7 0.035 2.7 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.7 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 2.195 1.115 2.195 0.93 2.125 0.93 2.125 1.065 1.915 1.065 1.915 0.925 1.78 0.925 1.78 0.825 1.31 0.825 1.31 0.475 1.655 0.475 1.655 0.29 1.585 0.29 1.585 0.425 1.375 0.425 1.375 0.36 1.325 0.36 1.325 0.425 1.26 0.425 1.26 0.875 1.73 0.875 1.73 0.975 1.865 0.975 1.865 1.115 ;
      POLYGON 1.655 1.105 1.655 0.925 1.105 0.925 1.105 0.725 0.63 0.725 0.63 0.475 0.835 0.475 0.835 0.375 1.105 0.375 1.105 0.3 1.375 0.3 1.375 0.135 1.865 0.135 1.865 0.26 1.915 0.26 1.915 0.135 2.125 0.135 2.125 0.275 2.195 0.275 2.195 0.085 1.325 0.085 1.325 0.25 1.105 0.25 1.105 0.185 1.055 0.185 1.055 0.325 0.835 0.325 0.835 0.275 0.785 0.275 0.785 0.425 0.58 0.425 0.58 0.525 0.15 0.525 0.15 0.575 0.58 0.575 0.58 0.775 0.785 0.775 0.785 0.9 0.835 0.9 0.835 0.775 1.055 0.775 1.055 0.975 1.325 0.975 1.325 1.1 1.375 1.1 1.375 0.975 1.585 0.975 1.585 1.105 ;
      POLYGON 0.565 1.015 0.565 0.825 0.09 0.825 0.09 0.375 0.565 0.375 0.565 0.185 0.515 0.185 0.515 0.325 0.295 0.325 0.295 0.2 0.245 0.2 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1 0.295 1 0.295 0.875 0.515 0.875 0.515 1.015 ;
      POLYGON 2.455 0.965 2.455 0.805 2.62 0.805 2.62 0.375 2.455 0.375 2.455 0.195 2.405 0.195 2.405 0.425 2.57 0.425 2.57 0.755 2.405 0.755 2.405 0.965 ;
      RECT 1.375 0.525 1.73 0.595 ;
    LAYER M2 ;
      RECT 0.335 0.825 1.49 0.875 ;
      RECT 1.5 0.525 2.66 0.575 ;
    LAYER VIA1 ;
      RECT 1.31 0.825 1.44 0.875 ;
      RECT 0.385 0.825 0.515 0.875 ;
      RECT 2.57 0.525 2.62 0.575 ;
      RECT 1.55 0.525 1.68 0.575 ;
  END
END XOR2_X4M_A12TL_C35

MACRO INV_X0P5B_A12TH_C35
  CLASS CORE ;
  FOREIGN INV_X0P5B_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.07 0.295 0.925 0.365 0.925 0.365 0.09 0.23 0.09 0.23 0.17 0.31 0.17 0.31 0.875 0.245 0.875 0.245 1.07 ;
    END
    ANTENNADIFFAREA 0.028125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.885 0.1 0.885 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.175 0.165 0.175 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.095 0.035 0.095 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P5B_A12TH_C35

MACRO INV_X6M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X6M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.5 0.525 0.5 0.425 0.28 0.425 0.28 0.475 0.45 0.475 0.45 0.525 0.145 0.525 0.145 0.575 0.72 0.575 0.72 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1932 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.01 0.295 0.875 0.515 0.875 0.515 0.995 0.565 0.995 0.565 0.875 0.785 0.875 0.785 0.995 0.835 0.995 0.835 0.875 1.04 0.875 1.04 0.32 0.835 0.32 0.835 0.2 0.785 0.2 0.785 0.32 0.565 0.32 0.565 0.2 0.515 0.2 0.515 0.32 0.295 0.32 0.295 0.185 0.245 0.185 0.245 0.375 0.985 0.375 0.985 0.82 0.245 0.82 0.245 1.01 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
END INV_X6M_A12TL_C35

MACRO INV_X5M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.161 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.85 0.375 0.85 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
END INV_X5M_A12TL_C35

MACRO INV_X7P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X7P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.675 1.04 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.77 0.525 0.77 0.425 0.55 0.425 0.55 0.475 0.72 0.475 0.72 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2422 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1 0.295 0.88 0.515 0.88 0.515 0.985 0.565 0.985 0.565 0.88 0.785 0.88 0.785 0.985 0.835 0.985 0.835 0.88 1.055 0.88 1.055 0.985 1.105 0.985 1.105 0.88 1.325 0.88 1.325 0.305 1.105 0.305 1.105 0.2 1.055 0.2 1.055 0.305 0.835 0.305 0.835 0.2 0.785 0.2 0.785 0.305 0.565 0.305 0.565 0.2 0.515 0.2 0.515 0.305 0.295 0.305 0.295 0.185 0.245 0.185 0.245 0.375 1.255 0.375 1.255 0.81 0.245 0.81 0.245 1 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.245 0.44 0.245 0.44 0.035 0.64 0.035 0.64 0.245 0.71 0.245 0.71 0.035 0.91 0.035 0.91 0.245 0.98 0.245 0.98 0.035 1.175 0.035 1.175 0.255 1.255 0.255 1.255 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
END INV_X7P5M_A12TL_C35

MACRO INV_X4B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X4B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.144 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.275 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.275 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X4B_A12TUL_C35

MACRO INV_X3P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X3P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.155 0.515 0.155 0.515 0.325 0.295 0.325 0.295 0.155 0.245 0.155 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.126 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.265 0.44 0.035 0.64 0.035 0.64 0.21 0.71 0.21 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.37 0.035 0.37 0.265 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X3P5B_A12TUL_C35

MACRO NOR2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.38 0.635 0.38 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.325 0.295 0.325 0.295 0.105 0.245 0.105 0.245 0.375 0.445 0.375 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.06025 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X1M_A12TUL_C35

MACRO OAI22_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.8 0.605 0.8 0.525 0.635 0.525 0.635 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.705 1.04 0.475 1.39 0.475 1.39 0.575 1.61 0.575 1.61 0.495 1.445 0.495 1.445 0.425 0.985 0.425 0.985 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.715 0.675 1.715 0.49 1.66 0.49 1.66 0.625 1.325 0.625 1.325 0.525 1.09 0.525 1.09 0.605 1.255 0.605 1.255 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.92 0.875 0.92 1 0.97 1 0.97 0.875 1.46 0.875 1.46 1 1.51 1 1.51 0.875 1.85 0.875 1.85 0.325 1.645 0.325 1.645 0.2 1.595 0.2 1.595 0.325 1.375 0.325 1.375 0.2 1.325 0.2 1.325 0.325 1.115 0.325 1.115 0.195 1.045 0.195 1.045 0.375 1.795 0.375 1.795 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.261 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.79 1.165 1.79 0.925 1.72 0.925 1.72 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.775 0.1 0.775 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.255 0.845 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.97 0.375 0.97 0.135 1.19 0.135 1.19 0.26 1.24 0.26 1.24 0.135 1.46 0.135 1.46 0.26 1.51 0.26 1.51 0.135 1.72 0.135 1.72 0.275 1.79 0.275 1.79 0.085 0.92 0.085 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OAI22_X3M_A12TUL_C35

MACRO OAI22_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.07 0.675 1.07 0.525 0.87 0.525 0.87 0.475 1.04 0.475 1.04 0.425 0.82 0.425 0.82 0.575 1.02 0.575 1.02 0.625 0.955 0.625 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.775 1.175 0.495 1.12 0.495 1.12 0.725 0.77 0.725 0.77 0.495 0.715 0.495 0.715 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.92 0.875 0.92 1 0.97 1 0.97 0.875 1.31 0.875 1.31 0.325 1.105 0.325 1.105 0.2 1.055 0.2 1.055 0.325 0.845 0.325 0.845 0.195 0.775 0.195 0.775 0.375 1.255 0.375 1.255 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.174 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 0.375 0.7 0.135 0.92 0.135 0.92 0.26 0.97 0.26 0.97 0.135 1.18 0.135 1.18 0.275 1.25 0.275 1.25 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OAI22_X2M_A12TUL_C35

MACRO AO21A1AI2_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.8 0.605 0.8 0.525 0.635 0.525 0.635 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.625 1.005 0.625 1.005 0.575 1.34 0.575 1.34 0.425 1.225 0.425 1.225 0.475 1.29 0.475 1.29 0.525 0.955 0.525 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.745 0.775 1.745 0.705 1.45 0.705 1.45 0.595 1.745 0.595 1.745 0.525 1.39 0.525 1.39 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.645 1.015 1.645 0.875 1.85 0.875 1.85 0.325 1.78 0.325 1.78 0.2 1.73 0.2 1.73 0.325 1.52 0.325 1.52 0.19 1.45 0.19 1.45 0.375 1.795 0.375 1.795 0.825 1.045 0.825 1.045 1.01 1.115 1.01 1.115 0.875 1.325 0.875 1.325 1 1.375 1 1.375 0.875 1.595 0.875 1.595 1.015 ;
    END
    ANTENNADIFFAREA 0.19975 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.79 1.165 1.79 0.93 1.72 0.93 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 1.25 0.255 1.25 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.115 1.25 0.93 1.18 0.93 1.18 1.065 0.97 1.065 0.97 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.115 ;
      POLYGON 1.375 0.375 1.375 0.135 1.585 0.135 1.585 0.27 1.655 0.27 1.655 0.085 1.325 0.085 1.325 0.325 1.105 0.325 1.105 0.2 1.055 0.2 1.055 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END AO21A1AI2_X3M_A12TUL_C35

MACRO INV_X7P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X7P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.675 1.04 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.77 0.525 0.77 0.425 0.55 0.425 0.55 0.475 0.72 0.475 0.72 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1904 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.31 0.875 1.31 0.325 1.105 0.325 1.105 0.095 1.055 0.095 1.055 0.325 0.835 0.325 0.835 0.095 0.785 0.095 0.785 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 1.255 0.375 1.255 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.272 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.22 1.25 0.22 1.25 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.22 0.17 0.22 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
END INV_X7P5B_A12TUL_C35

MACRO AOI21_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.8 0.605 0.8 0.525 0.635 0.525 0.635 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.625 1.005 0.625 1.005 0.575 1.34 0.575 1.34 0.425 1.225 0.425 1.225 0.475 1.29 0.475 1.29 0.525 0.955 0.525 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.07665 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.115 1.005 1.115 0.875 1.325 0.875 1.325 1 1.375 1 1.375 0.875 1.445 0.875 1.445 0.325 1.24 0.325 1.24 0.105 1.19 0.105 1.19 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 1.39 0.375 1.39 0.825 1.045 0.825 1.045 1.005 ;
    END
    ANTENNADIFFAREA 0.17975 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.315 0.035 1.315 0.27 1.385 0.27 1.385 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.115 1.25 0.935 1.18 0.935 1.18 1.065 0.97 1.065 0.97 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.115 ;
  END
END AOI21_X3M_A12TUL_C35

MACRO OAI22_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.43 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.605 1.07 0.605 1.07 0.525 0.835 0.525 0.835 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1218 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.705 1.175 0.425 0.715 0.425 0.715 0.555 0.635 0.555 0.635 0.425 0.175 0.425 0.175 0.705 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.77 0.605 0.77 0.475 1.12 0.475 1.12 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1218 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.985 0.675 1.985 0.605 2.15 0.605 2.15 0.525 1.915 0.525 1.915 0.625 1.595 0.625 1.595 0.525 1.36 0.525 1.36 0.605 1.525 0.605 1.525 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1218 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.255 0.705 2.255 0.425 1.795 0.425 1.795 0.525 1.715 0.525 1.715 0.425 1.255 0.425 1.255 0.705 1.31 0.705 1.31 0.475 1.66 0.475 1.66 0.575 1.85 0.575 1.85 0.475 2.2 0.475 2.2 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1218 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.92 0.875 0.92 1 0.97 1 0.97 0.875 1.46 0.875 1.46 1 1.51 1 1.51 0.875 2 0.875 2 1 2.05 1 2.05 0.875 2.39 0.875 2.39 0.325 2.185 0.325 2.185 0.2 2.135 0.2 2.135 0.325 1.915 0.325 1.915 0.2 1.865 0.2 1.865 0.325 1.645 0.325 1.645 0.2 1.595 0.2 1.595 0.325 1.385 0.325 1.385 0.195 1.315 0.195 1.315 0.375 2.335 0.375 2.335 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.348 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
      LAYER M1 ;
        POLYGON 2.43 1.235 2.43 1.165 2.33 1.165 2.33 0.93 2.26 0.93 2.26 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.775 0.1 0.775 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.43 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
      LAYER M1 ;
        POLYGON 1.115 0.255 1.115 0.035 2.43 0.035 2.43 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 2.43 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.24 0.375 1.24 0.135 1.46 0.135 1.46 0.26 1.51 0.26 1.51 0.135 1.73 0.135 1.73 0.26 1.78 0.26 1.78 0.135 2 0.135 2 0.26 2.05 0.26 2.05 0.135 2.26 0.135 2.26 0.27 2.33 0.27 2.33 0.085 1.19 0.085 1.19 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OAI22_X4M_A12TUL_C35

MACRO INV_X6B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X6B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.5 0.525 0.5 0.425 0.28 0.425 0.28 0.475 0.45 0.475 0.45 0.525 0.145 0.525 0.145 0.575 0.72 0.575 0.72 0.625 0.55 0.625 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1512 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.095 0.785 0.095 0.785 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.985 0.375 0.985 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.275 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.275 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
END INV_X6B_A12TUL_C35

MACRO XOR2_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.295 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.67 0.625 1.8 0.675 ;
        RECT 2.055 0.625 2.105 0.675 ;
      LAYER M1 ;
        POLYGON 1.85 0.675 1.85 0.485 1.8 0.485 1.8 0.625 1.58 0.625 1.58 0.485 1.53 0.485 1.53 0.675 ;
        RECT 2.045 0.435 2.115 0.725 ;
      LAYER M2 ;
        RECT 1.62 0.625 2.16 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 LAYER M1 ;
    ANTENNAGATEAREA 0.09625 LAYER M2 ;
    ANTENNAGATEAREA 0.09625 LAYER M3 ;
    ANTENNAGATEAREA 0.09625 LAYER M4 ;
    ANTENNAGATEAREA 0.09625 LAYER M5 ;
    ANTENNAGATEAREA 0.09625 LAYER M6 ;
    ANTENNAGATEAREA 0.09625 LAYER M7 ;
    ANTENNAGATEAREA 0.09625 LAYER M8 ;
    ANTENNAGATEAREA 0.09625 LAYER AP ;
    ANTENNAMAXAREACAR 0.6304348 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2018634 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.675 0.77 0.625 0.6 0.625 0.6 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.55 0.525 0.55 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.78 1 1.78 0.875 1.985 0.875 1.985 0.325 1.78 0.325 1.78 0.2 1.73 0.2 1.73 0.325 1.51 0.325 1.51 0.185 1.18 0.185 1.18 0.365 1.25 0.365 1.25 0.235 1.46 0.235 1.46 0.375 1.93 0.375 1.93 0.825 1.16 0.825 1.16 0.875 1.73 0.875 1.73 1 ;
    END
    ANTENNADIFFAREA 0.183 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
      LAYER M1 ;
        POLYGON 2.295 1.235 2.295 1.165 2.06 1.165 2.06 0.93 1.99 0.93 1.99 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.295 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.335 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.99 0.035 1.99 0.275 2.06 0.275 2.06 0.035 2.295 0.035 2.295 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 2.295 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.93 1.115 1.93 0.925 1.85 0.925 1.85 1.065 1.645 1.065 1.645 0.925 1.07 0.925 1.07 0.475 1.385 0.475 1.385 0.295 1.315 0.295 1.315 0.425 1.115 0.425 1.115 0.185 1.045 0.185 1.045 0.425 1.02 0.425 1.02 0.975 1.595 0.975 1.595 1.115 ;
      POLYGON 1.405 1.075 1.405 1.025 0.97 1.025 0.97 0.825 0.565 0.825 0.565 0.725 0.495 0.725 0.495 0.455 0.7 0.455 0.7 0.375 0.97 0.375 0.97 0.135 1.595 0.135 1.595 0.26 1.645 0.26 1.645 0.135 1.855 0.135 1.855 0.275 1.925 0.275 1.925 0.085 0.92 0.085 0.92 0.325 0.7 0.325 0.7 0.265 0.65 0.265 0.65 0.405 0.445 0.405 0.445 0.525 0.15 0.525 0.15 0.575 0.445 0.575 0.445 0.775 0.515 0.775 0.515 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.075 ;
      POLYGON 0.43 1.025 0.43 0.825 0.09 0.825 0.09 0.355 0.43 0.355 0.43 0.165 0.38 0.165 0.38 0.305 0.16 0.305 0.16 0.18 0.11 0.18 0.11 0.305 0.04 0.305 0.04 0.875 0.11 0.875 0.11 1.025 0.16 1.025 0.16 0.875 0.38 0.875 0.38 1.025 ;
      POLYGON 2.185 0.985 2.185 0.845 2.215 0.845 2.215 0.315 2.185 0.315 2.185 0.175 2.135 0.175 2.135 0.365 2.165 0.365 2.165 0.795 2.135 0.795 2.135 0.985 ;
      POLYGON 1.445 0.715 1.445 0.525 1.125 0.525 1.125 0.715 1.175 0.715 1.175 0.575 1.395 0.575 1.395 0.715 ;
    LAYER M2 ;
      RECT 0.06 0.925 1.25 0.975 ;
      RECT 1.215 0.525 2.255 0.575 ;
    LAYER VIA1 ;
      RECT 1.07 0.925 1.2 0.975 ;
      RECT 0.38 0.925 0.43 0.975 ;
      RECT 0.11 0.925 0.16 0.975 ;
      RECT 2.165 0.525 2.215 0.575 ;
      RECT 1.265 0.525 1.395 0.575 ;
  END
END XOR2_X3M_A12TUL_C35

MACRO OA21A1OI2_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.8 0.605 0.8 0.525 0.635 0.525 0.635 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.625 1.005 0.625 1.005 0.575 1.34 0.575 1.34 0.425 1.225 0.425 1.225 0.475 1.29 0.475 1.29 0.525 0.955 0.525 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.58 0.675 1.58 0.575 1.745 0.575 1.745 0.425 1.63 0.425 1.63 0.475 1.695 0.475 1.695 0.525 1.455 0.525 1.455 0.485 1.39 0.485 1.39 0.575 1.53 0.575 1.53 0.625 1.36 0.625 1.36 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.07665 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.52 1.005 1.52 0.875 1.73 0.875 1.73 1 1.78 1 1.78 0.875 1.85 0.875 1.85 0.325 1.645 0.325 1.645 0.185 1.595 0.185 1.595 0.325 1.375 0.325 1.375 0.2 1.325 0.2 1.325 0.325 1.115 0.325 1.115 0.195 1.045 0.195 1.045 0.375 1.795 0.375 1.795 0.825 1.45 0.825 1.45 1.005 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 1.79 0.27 1.79 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.45 0.035 1.45 0.27 1.52 0.27 1.52 0.035 1.72 0.035 1.72 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.655 1.11 1.655 0.93 1.585 0.93 1.585 1.06 1.375 1.06 1.375 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.325 0.875 1.325 1.11 ;
      POLYGON 0.97 0.375 0.97 0.14 1.18 0.14 1.18 0.275 1.25 0.275 1.25 0.09 0.92 0.09 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OA21A1OI2_X3M_A12TUL_C35

MACRO NAND2_X2A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X2A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.77 0.875 0.77 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.103 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X2A_A12TUL_C35

MACRO OAI22_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI22_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.07 0.675 1.07 0.525 0.87 0.525 0.87 0.475 1.04 0.475 1.04 0.425 0.82 0.425 0.82 0.575 1.02 0.575 1.02 0.625 0.955 0.625 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.775 1.175 0.495 1.12 0.495 1.12 0.725 0.77 0.725 0.77 0.495 0.715 0.495 0.715 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.92 0.875 0.92 1 0.97 1 0.97 0.875 1.31 0.875 1.31 0.325 1.105 0.325 1.105 0.225 1.055 0.225 1.055 0.325 0.835 0.325 0.835 0.225 0.785 0.225 0.785 0.375 1.255 0.375 1.255 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.25 1.165 1.25 0.93 1.18 0.93 1.18 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 0.375 0.7 0.135 0.92 0.135 0.92 0.26 0.97 0.26 0.97 0.135 1.18 0.135 1.18 0.27 1.25 0.27 1.25 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.14 0.38 0.14 0.38 0.325 0.16 0.325 0.16 0.13 0.11 0.13 0.11 0.375 ;
  END
END OAI22_X1P4M_A12TUL_C35

MACRO AOI21_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI21_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.675 0.905 0.625 0.735 0.625 0.735 0.575 0.935 0.575 0.935 0.425 0.82 0.425 0.82 0.475 0.885 0.475 0.885 0.525 0.685 0.525 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0511 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.105 0.785 0.105 0.785 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.985 0.375 0.985 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.109 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.98 1.115 0.98 0.93 0.91 0.93 0.91 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
  END
END AOI21_X2M_A12TUL_C35

MACRO XOR2_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.185 0.625 0.235 0.675 ;
        RECT 1.285 0.625 1.415 0.675 ;
      LAYER M1 ;
        POLYGON 1.455 0.675 1.455 0.485 1.395 0.485 1.395 0.625 1.305 0.625 1.305 0.485 1.245 0.485 1.245 0.675 ;
        RECT 0.18 0.425 0.24 0.725 ;
      LAYER M2 ;
        RECT 0.135 0.625 1.465 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 LAYER M1 ;
    ANTENNAGATEAREA 0.0763 LAYER M2 ;
    ANTENNAGATEAREA 0.0763 LAYER M3 ;
    ANTENNAGATEAREA 0.0763 LAYER M4 ;
    ANTENNAGATEAREA 0.0763 LAYER M5 ;
    ANTENNAGATEAREA 0.0763 LAYER M6 ;
    ANTENNAGATEAREA 0.0763 LAYER M7 ;
    ANTENNAGATEAREA 0.0763 LAYER M8 ;
    ANTENNAGATEAREA 0.0763 LAYER AP ;
    ANTENNAMAXAREACAR 0.612245 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2210884 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.805 0.365 0.595 0.53 0.595 0.53 0.525 0.295 0.525 0.295 0.595 0.31 0.595 0.31 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.51 1.105 1.51 0.905 1.58 0.905 1.58 0.295 1.51 0.295 1.51 0.115 0.985 0.115 0.985 0.085 0.905 0.085 0.905 0.165 1.46 0.165 1.46 0.345 1.525 0.345 1.525 0.855 1.46 0.855 1.46 1.055 1.24 1.055 1.24 0.93 1.19 0.93 1.19 1.055 0.985 1.055 0.985 1.025 0.905 1.025 0.905 1.105 ;
    END
    ANTENNADIFFAREA 0.1675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 0.85 1.165 0.85 1.03 0.77 1.03 0.77 1.165 0.575 1.165 0.575 1.045 0.505 1.045 0.505 1.165 0.305 1.165 0.305 0.875 0.235 0.875 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.16 0.575 0.16 0.575 0.035 0.77 0.035 0.77 0.17 0.85 0.17 0.85 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 1.105 0.44 0.975 1.04 0.975 1.04 1 1.12 1 1.12 0.83 1.04 0.83 1.04 0.925 0.55 0.925 0.55 0.725 0.635 0.725 0.635 0.585 0.785 0.585 0.785 0.515 0.635 0.515 0.635 0.425 0.43 0.425 0.43 0.275 1.315 0.275 1.315 0.405 1.385 0.405 1.385 0.225 0.38 0.225 0.38 0.475 0.585 0.475 0.585 0.675 0.5 0.675 0.5 0.925 0.37 0.925 0.37 1.105 ;
      POLYGON 0.16 0.985 0.16 0.795 0.13 0.795 0.13 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.08 0.305 0.08 0.845 0.11 0.845 0.11 0.985 ;
      POLYGON 1.375 0.975 1.375 0.725 0.9 0.725 0.9 0.375 1.135 0.375 1.135 0.325 0.62 0.325 0.62 0.375 0.85 0.375 0.85 0.805 0.62 0.805 0.62 0.855 0.9 0.855 0.9 0.775 1.325 0.775 1.325 0.975 ;
      POLYGON 1.185 0.625 1.185 0.425 0.975 0.425 0.975 0.625 1.035 0.625 1.035 0.475 1.125 0.475 1.125 0.625 ;
    LAYER M2 ;
      RECT 0.04 0.425 1.195 0.475 ;
    LAYER VIA1 ;
      RECT 1.015 0.425 1.145 0.475 ;
      RECT 0.08 0.425 0.13 0.475 ;
  END
END XOR2_X2M_A12TUL_C35

MACRO INV_X16M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X16M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.12 0.675 2.12 0.58 2.18 0.58 2.18 0.6 2.27 0.6 2.27 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 0.5 0.675 0.5 0.575 0.99 0.575 0.99 0.625 0.82 0.625 0.82 0.675 1.04 0.675 1.04 0.575 1.53 0.575 1.53 0.625 1.36 0.625 1.36 0.675 1.58 0.675 1.58 0.575 2.07 0.575 2.07 0.625 1.9 0.625 1.9 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5152 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 0.935 0.295 0.885 0.515 0.885 0.515 0.93 0.565 0.93 0.565 0.885 0.785 0.885 0.785 0.93 0.835 0.93 0.835 0.885 1.055 0.885 1.055 0.93 1.105 0.93 1.105 0.885 1.325 0.885 1.325 0.93 1.375 0.93 1.375 0.885 1.595 0.885 1.595 0.93 1.645 0.93 1.645 0.885 1.865 0.885 1.865 0.93 1.915 0.93 1.915 0.885 2.135 0.885 2.135 0.93 2.185 0.93 2.185 0.885 2.46 0.885 2.46 0.315 2.185 0.315 2.185 0.27 2.135 0.27 2.135 0.315 1.915 0.315 1.915 0.27 1.865 0.27 1.865 0.315 1.645 0.315 1.645 0.27 1.595 0.27 1.595 0.315 1.375 0.315 1.375 0.27 1.325 0.27 1.325 0.315 1.105 0.315 1.105 0.27 1.055 0.27 1.055 0.315 0.835 0.315 0.835 0.27 0.785 0.27 0.785 0.315 0.565 0.315 0.565 0.27 0.515 0.27 0.515 0.315 0.295 0.315 0.295 0.265 0.245 0.265 0.245 0.455 2.325 0.455 2.325 0.745 0.245 0.745 0.245 0.935 ;
    END
    ANTENNADIFFAREA 0.736 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
      LAYER M1 ;
        POLYGON 2.565 1.235 2.565 1.165 2.465 1.165 2.465 0.995 2.395 0.995 2.395 1.165 2.33 1.165 2.33 0.945 2.26 0.945 2.26 1.165 2.06 1.165 2.06 0.945 1.99 0.945 1.99 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.565 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 1.72 0.035 1.72 0.255 1.79 0.255 1.79 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.26 0.035 2.26 0.255 2.33 0.255 2.33 0.035 2.395 0.035 2.395 0.205 2.465 0.205 2.465 0.035 2.565 0.035 2.565 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 2.565 0.065 ;
    END
  END VSS
END INV_X16M_A12TUL_C35

MACRO INV_X3B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X3B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.575 0.325 0.575 0.09 0.505 0.09 0.505 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.126 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X3B_A12TUL_C35

MACRO INV_X5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.845 0.325 0.845 0.09 0.775 0.09 0.775 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.85 0.375 0.85 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.198 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.275 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.275 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
END INV_X5B_A12TUL_C35

MACRO NAND2_X1P4B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1P4B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.425 0.28 0.425 0.28 0.495 0.445 0.495 0.445 0.605 0.28 0.605 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0427 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0427 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.093 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.94 0.37 0.94 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X1P4B_A12TUL_C35

MACRO INV_X13M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X13M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.16 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.715 0.675 1.715 0.58 1.86 0.58 1.86 0.5 1.78 0.5 1.78 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 0.635 0.675 0.635 0.575 1.125 0.575 1.125 0.625 0.955 0.625 0.955 0.675 1.175 0.675 1.175 0.575 1.665 0.575 1.665 0.625 1.495 0.625 1.495 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4186 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 0.96 0.295 0.885 0.515 0.885 0.515 0.95 0.565 0.95 0.565 0.885 0.785 0.885 0.785 0.95 0.835 0.95 0.835 0.885 1.055 0.885 1.055 0.95 1.105 0.95 1.105 0.885 1.325 0.885 1.325 0.95 1.375 0.95 1.375 0.885 1.595 0.885 1.595 0.95 1.645 0.95 1.645 0.885 1.865 0.885 1.865 0.95 1.915 0.95 1.915 0.885 2.05 0.885 2.05 0.285 2 0.285 2 0.315 1.915 0.315 1.915 0.25 1.865 0.25 1.865 0.315 1.645 0.315 1.645 0.25 1.595 0.25 1.595 0.315 1.375 0.315 1.375 0.25 1.325 0.25 1.325 0.315 1.105 0.315 1.105 0.25 1.055 0.25 1.055 0.315 0.835 0.315 0.835 0.25 0.785 0.25 0.785 0.315 0.565 0.315 0.565 0.25 0.515 0.25 0.515 0.315 0.295 0.315 0.295 0.215 0.245 0.215 0.245 0.43 1.93 0.43 1.93 0.77 0.245 0.77 0.245 0.96 ;
    END
    ANTENNADIFFAREA 0.713 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
      LAYER M1 ;
        POLYGON 2.16 1.235 2.16 1.165 1.79 1.165 1.79 0.945 1.72 0.945 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.16 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 1.72 0.035 1.72 0.255 1.79 0.255 1.79 0.035 2.16 0.035 2.16 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 2.16 0.065 ;
    END
  END VSS
END INV_X13M_A12TUL_C35

MACRO INV_X1P4B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P4B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.225 0.295 0.225 0.295 0.11 0.245 0.11 0.245 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.051 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.195 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P4B_A12TUL_C35

MACRO INV_X1P7B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P7B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.605 0.145 0.605 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04235 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.225 0.295 0.225 0.295 0.145 0.245 0.145 0.245 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.0605 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.205 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.205 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P7B_A12TUL_C35

MACRO INV_X2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.095 0.245 0.095 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.072 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X2B_A12TUL_C35

MACRO NAND2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0238 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0238 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.04 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.825 0.245 0.825 0.245 1.04 ;
    END
    ANTENNADIFFAREA 0.05775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.87 0.1 0.87 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X1M_A12TUL_C35

MACRO INV_X2P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X2P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.565 0.325 0.565 0.135 0.515 0.135 0.515 0.325 0.295 0.325 0.295 0.145 0.245 0.145 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.2 0.17 0.2 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X2P5B_A12TUL_C35

MACRO INV_X1P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05425 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.0775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P7M_A12TUL_C35

MACRO AO21B_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.725 0.33 0.725 0.33 0.675 0.53 0.675 0.53 0.525 0.415 0.525 0.415 0.575 0.48 0.575 0.48 0.625 0.28 0.625 0.28 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05145 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.65 0.605 0.65 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05145 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.61 0.605 1.61 0.525 1.445 0.525 1.445 0.425 0.985 0.425 0.985 0.525 0.82 0.525 0.82 0.605 1.04 0.605 1.04 0.475 1.39 0.475 1.39 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1204 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.015 0.835 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.325 0.875 1.325 1 1.375 1 1.375 0.875 1.595 0.875 1.595 1 1.645 1 1.645 0.875 1.85 0.875 1.85 0.325 1.51 0.325 1.51 0.2 1.46 0.2 1.46 0.325 0.97 0.325 0.97 0.185 0.92 0.185 0.92 0.375 1.795 0.375 1.795 0.825 0.785 0.825 0.785 1.015 ;
    END
    ANTENNADIFFAREA 0.262 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 1.79 1.165 1.79 0.93 1.72 0.93 1.72 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.355 0.71 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.72 0.035 1.72 0.27 1.79 0.27 1.79 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.64 0.035 0.64 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1 0.565 0.875 0.7 0.875 0.7 0.725 1.17 0.725 1.17 0.615 1.255 0.615 1.255 0.725 1.71 0.725 1.71 0.565 1.66 0.565 1.66 0.675 1.305 0.675 1.305 0.565 1.12 0.565 1.12 0.675 0.765 0.675 0.765 0.565 0.715 0.565 0.715 0.675 0.65 0.675 0.65 0.825 0.09 0.825 0.09 0.375 0.43 0.375 0.43 0.185 0.38 0.185 0.38 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1 0.295 1 0.295 0.875 0.515 0.875 0.515 1 ;
  END
END AO21B_X4M_A12TUL_C35

MACRO XOR2_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR2_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.62 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.19 0.625 0.24 0.675 ;
        RECT 1.285 0.625 1.415 0.675 ;
      LAYER M1 ;
        POLYGON 1.455 0.675 1.455 0.485 1.395 0.485 1.395 0.625 1.305 0.625 1.305 0.485 1.245 0.485 1.245 0.675 ;
        RECT 0.18 0.425 0.25 0.725 ;
      LAYER M2 ;
        RECT 0.14 0.625 1.47 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02905 LAYER M1 ;
    ANTENNAGATEAREA 0.0651 LAYER M2 ;
    ANTENNAGATEAREA 0.0651 LAYER M3 ;
    ANTENNAGATEAREA 0.0651 LAYER M4 ;
    ANTENNAGATEAREA 0.0651 LAYER M5 ;
    ANTENNAGATEAREA 0.0651 LAYER M6 ;
    ANTENNAGATEAREA 0.0651 LAYER M7 ;
    ANTENNAGATEAREA 0.0651 LAYER M8 ;
    ANTENNAGATEAREA 0.0651 LAYER AP ;
    ANTENNAMAXAREACAR 0.7572815 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2237522 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.805 0.365 0.575 0.53 0.575 0.53 0.525 0.31 0.525 0.31 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04515 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.51 1.105 1.51 0.905 1.58 0.905 1.58 0.295 1.51 0.295 1.51 0.11 0.99 0.11 0.99 0.09 0.9 0.09 0.9 0.16 1.46 0.16 1.46 0.345 1.525 0.345 1.525 0.855 1.46 0.855 1.46 1.055 1.24 1.055 1.24 0.93 1.19 0.93 1.19 1.055 0.985 1.055 0.985 1.025 0.905 1.025 0.905 1.105 ;
    END
    ANTENNADIFFAREA 0.13425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
      LAYER M1 ;
        POLYGON 1.62 1.235 1.62 1.165 0.85 1.165 0.85 1.03 0.77 1.03 0.77 1.165 0.575 1.165 0.575 1.045 0.505 1.045 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.62 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.5 0.035 0.5 0.155 0.58 0.155 0.58 0.035 0.77 0.035 0.77 0.155 0.85 0.155 0.85 0.035 1.62 0.035 1.62 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.62 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 1.105 0.44 0.975 1.04 0.975 1.04 1 1.12 1 1.12 0.83 1.04 0.83 1.04 0.925 0.55 0.925 0.55 0.695 0.765 0.695 0.765 0.425 0.43 0.425 0.43 0.26 1.325 0.26 1.325 0.4 1.375 0.4 1.375 0.21 0.43 0.21 0.43 0.165 0.38 0.165 0.38 0.475 0.715 0.475 0.715 0.645 0.5 0.645 0.5 0.925 0.37 0.925 0.37 1.105 ;
      POLYGON 1.39 0.995 1.39 0.83 1.36 0.83 1.36 0.725 0.9 0.725 0.9 0.36 1.135 0.36 1.135 0.31 0.62 0.31 0.62 0.36 0.85 0.36 0.85 0.805 0.62 0.805 0.62 0.855 0.9 0.855 0.9 0.775 1.31 0.775 1.31 0.995 ;
      POLYGON 0.16 0.985 0.16 0.795 0.13 0.795 0.13 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.08 0.305 0.08 0.845 0.11 0.845 0.11 0.985 ;
      POLYGON 1.185 0.615 1.185 0.425 0.975 0.425 0.975 0.615 1.035 0.615 1.035 0.475 1.125 0.475 1.125 0.615 ;
    LAYER M2 ;
      RECT 0.04 0.425 1.195 0.475 ;
    LAYER VIA1 ;
      RECT 1.015 0.425 1.145 0.475 ;
      RECT 0.08 0.425 0.13 0.475 ;
  END
END XOR2_X1P4M_A12TUL_C35

MACRO INV_X1B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0252 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.225 0.305 0.225 0.305 0.09 0.235 0.09 0.235 0.275 0.31 0.275 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.054 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X1B_A12TUL_C35

MACRO AO1B2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO1B2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0147 ;
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 0.975 0.77 0.975 0.77 0.295 0.7 0.295 0.7 0.155 0.65 0.155 0.65 0.345 0.715 0.345 0.715 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.07575 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.095 0.295 0.875 0.63 0.875 0.63 0.565 0.58 0.565 0.58 0.825 0.075 0.825 0.075 0.24 0.19 0.24 0.19 0.19 0.025 0.19 0.025 0.875 0.245 0.875 0.245 1.095 ;
  END
END AO1B2_X1M_A12TUL_C35

MACRO INV_X1P2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.225 0.295 0.225 0.295 0.095 0.245 0.095 0.245 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.043 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.18 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P2B_A12TUL_C35

MACRO AOI22_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.07 0.675 1.07 0.525 0.87 0.525 0.87 0.475 1.04 0.475 1.04 0.425 0.82 0.425 0.82 0.575 1.02 0.575 1.02 0.625 0.955 0.625 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.775 1.175 0.495 1.12 0.495 1.12 0.725 0.77 0.725 0.77 0.495 0.715 0.495 0.715 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.31 0.875 1.31 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 1.255 0.375 1.255 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.174 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.42 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.18 0.035 1.18 0.27 1.25 0.27 1.25 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.42 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.115 1.25 0.925 1.18 0.925 1.18 1.065 0.97 1.065 0.97 0.94 0.92 0.94 0.92 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
  END
END AOI22_X2M_A12TUL_C35

MACRO BUFH_X7P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X7P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.575 0.8 0.575 0.8 0.425 0.685 0.425 0.685 0.475 0.75 0.475 0.75 0.525 0.365 0.525 0.365 0.425 0.145 0.425 0.145 0.475 0.315 0.475 0.315 0.525 0.145 0.525 0.145 0.575 0.585 0.575 0.585 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.139125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.97 0.995 0.97 0.875 1.19 0.875 1.19 0.98 1.24 0.98 1.24 0.875 1.46 0.875 1.46 0.98 1.51 0.98 1.51 0.875 1.73 0.875 1.73 0.98 1.78 0.98 1.78 0.875 1.99 0.875 1.99 0.325 1.78 0.325 1.78 0.22 1.73 0.22 1.73 0.325 1.51 0.325 1.51 0.22 1.46 0.22 1.46 0.325 1.24 0.325 1.24 0.22 1.19 0.22 1.19 0.325 0.97 0.325 0.97 0.205 0.92 0.205 0.92 0.395 1.92 0.395 1.92 0.805 0.92 0.805 0.92 0.995 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.925 1.165 1.925 0.93 1.855 0.93 1.855 1.165 1.655 1.165 1.655 0.945 1.585 0.945 1.585 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.945 1.045 0.945 1.045 1.165 0.845 1.165 0.845 0.845 0.775 0.845 0.775 1.165 0.575 1.165 0.575 0.845 0.505 0.845 0.505 1.165 0.305 1.165 0.305 0.845 0.235 0.845 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.355 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.585 0.035 1.585 0.255 1.655 0.255 1.655 0.035 1.855 0.035 1.855 0.27 1.925 0.27 1.925 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.7 0.9 0.7 0.775 0.835 0.775 0.835 0.675 0.9 0.675 0.9 0.585 1.785 0.585 1.785 0.625 1.855 0.625 1.855 0.535 0.85 0.535 0.85 0.625 0.785 0.625 0.785 0.725 0.075 0.725 0.075 0.375 0.7 0.375 0.7 0.185 0.65 0.185 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.2 0.11 0.2 0.11 0.325 0.025 0.325 0.025 0.775 0.11 0.775 0.11 0.9 0.16 0.9 0.16 0.775 0.38 0.775 0.38 0.9 0.43 0.9 0.43 0.775 0.65 0.775 0.65 0.9 ;
  END
END BUFH_X7P5M_A12TUL_C35

MACRO NAND2B_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2B_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.71 0.23 0.495 0.365 0.495 0.365 0.425 0.145 0.425 0.145 0.495 0.175 0.495 0.175 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.014525 ;
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.365 0.725 0.365 0.575 0.31 0.575 0.31 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0476 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.875 0.905 0.875 0.905 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.85 0.375 0.85 0.825 0.38 0.825 0.38 1.045 0.43 1.045 0.43 0.875 0.65 0.875 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.095 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.87 0.235 0.87 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.095 0.16 0.89 0.075 0.89 0.075 0.375 0.415 0.375 0.415 0.575 0.65 0.575 0.65 0.505 0.465 0.505 0.465 0.325 0.16 0.325 0.16 0.145 0.11 0.145 0.11 0.325 0.025 0.325 0.025 0.94 0.11 0.94 0.11 1.095 ;
  END
END NAND2B_X2M_A12TUL_C35

MACRO INV_X1P2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0385 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.13 0.245 0.13 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.055 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.305 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P2M_A12TUL_C35

MACRO INV_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0455 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.175 0.245 0.175 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P4M_A12TUL_C35

MACRO BUFH_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.525 0.145 0.525 0.145 0.575 0.345 0.575 0.345 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05565 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.85 0.375 0.85 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 0.705 0.565 0.705 0.605 0.775 0.605 0.775 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUFH_X3M_A12TUL_C35

MACRO AO21B_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.575 0.235 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.165 0.375 0.165 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.026075 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.445 0.31 0.445 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.026075 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.525 0.6 0.525 0.6 0.475 0.77 0.475 0.77 0.425 0.55 0.425 0.55 0.575 0.75 0.575 0.75 0.625 0.685 0.625 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0602 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.7 0.325 0.7 0.185 0.65 0.185 0.65 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.131 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.265 0.44 0.265 0.44 0.035 0.91 0.035 0.91 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1 0.295 0.875 0.465 0.875 0.465 0.775 0.9 0.775 0.9 0.565 0.85 0.565 0.85 0.725 0.495 0.725 0.495 0.565 0.445 0.565 0.445 0.725 0.415 0.725 0.415 0.825 0.075 0.825 0.075 0.275 0.17 0.275 0.17 0.095 0.1 0.095 0.1 0.225 0.025 0.225 0.025 0.875 0.245 0.875 0.245 1 ;
  END
END AO21B_X2M_A12TUL_C35

MACRO AOI22_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.425 0.28 0.425 0.28 0.495 0.445 0.495 0.445 0.605 0.28 0.605 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.675 1.04 0.425 0.82 0.425 0.82 0.495 0.985 0.495 0.985 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.775 1.175 0.495 1.12 0.495 1.12 0.725 0.77 0.725 0.77 0.495 0.715 0.495 0.715 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04305 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.005 0.845 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.31 0.875 1.31 0.325 0.97 0.325 0.97 0.14 0.92 0.14 0.92 0.325 0.43 0.325 0.43 0.14 0.38 0.14 0.38 0.375 1.255 0.375 1.255 0.825 0.775 0.825 0.775 1.005 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.315 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.18 0.035 1.18 0.27 1.25 0.27 1.25 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.315 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.25 1.115 1.25 0.925 1.18 0.925 1.18 1.065 0.97 1.065 0.97 0.94 0.92 0.94 0.92 1.065 0.7 1.065 0.7 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1.115 ;
  END
END AOI22_X1P4M_A12TUL_C35

MACRO XOR3_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XOR3_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.025 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.645 1.105 1.645 0.675 1.85 0.675 1.85 0.395 1.795 0.395 1.795 0.625 1.58 0.625 1.58 0.495 1.525 0.495 1.525 0.675 1.595 0.675 1.595 1.055 1.225 1.055 1.225 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.041475 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.805 0.23 0.575 0.65 0.575 0.65 0.505 0.56 0.505 0.56 0.52 0.175 0.52 0.175 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03955 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.85 0.495 0.85 0.605 0.82 0.605 0.82 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01925 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.525 0.995 1.525 0.825 1.31 0.825 1.31 0.375 1.405 0.375 1.405 0.325 1.255 0.325 1.255 0.875 1.45 0.875 1.45 0.995 ;
    END
    ANTENNADIFFAREA 0.068875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
      LAYER M1 ;
        POLYGON 2.025 1.235 2.025 1.165 1.79 1.165 1.79 0.845 1.72 0.845 1.72 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.875 0.235 0.875 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.025 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.345 0.305 0.035 0.905 0.035 0.905 0.17 0.985 0.17 0.985 0.035 1.72 0.035 1.72 0.29 1.79 0.29 1.79 0.035 2.025 0.035 2.025 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.345 ;
      LAYER M2 ;
        RECT 0 -0.065 2.025 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.115 1.105 1.115 0.975 1.305 0.975 1.305 0.995 1.395 0.995 1.395 0.925 1.17 0.925 1.17 0.275 1.49 0.275 1.49 0.425 1.66 0.425 1.66 0.505 1.71 0.505 1.71 0.375 1.54 0.375 1.54 0.225 1.24 0.225 1.24 0.1 1.19 0.1 1.19 0.22 1.115 0.22 1.115 0.09 1.045 0.09 1.045 0.27 1.12 0.27 1.12 0.925 1.045 0.925 1.045 1.105 ;
      POLYGON 0.43 1.085 0.43 0.945 0.565 0.945 0.565 0.755 0.515 0.755 0.515 0.895 0.38 0.895 0.38 1.085 ;
      POLYGON 0.16 1.075 0.16 0.885 0.105 0.885 0.105 0.465 0.43 0.465 0.43 0.135 0.795 0.135 0.795 0.085 0.38 0.085 0.38 0.415 0.16 0.415 0.16 0.25 0.11 0.25 0.11 0.415 0.055 0.415 0.055 0.935 0.11 0.935 0.11 1.075 ;
      POLYGON 0.7 1.015 0.7 0.875 1.04 0.875 1.04 0.325 0.985 0.325 0.985 0.225 0.515 0.225 0.515 0.415 0.565 0.415 0.565 0.275 0.935 0.275 0.935 0.375 0.99 0.375 0.99 0.825 0.65 0.825 0.65 1.015 ;
      POLYGON 1.915 0.935 1.915 0.775 1.985 0.775 1.985 0.175 1.85 0.175 1.85 0.255 1.935 0.255 1.935 0.725 1.755 0.725 1.755 0.775 1.865 0.775 1.865 0.935 ;
      POLYGON 1.525 0.775 1.525 0.725 1.45 0.725 1.45 0.47 1.38 0.47 1.38 0.775 ;
      POLYGON 0.865 0.775 0.865 0.725 0.76 0.725 0.76 0.375 0.865 0.375 0.865 0.325 0.63 0.325 0.63 0.395 0.71 0.395 0.71 0.635 0.285 0.635 0.285 0.705 0.395 0.705 0.395 0.685 0.71 0.685 0.71 0.775 ;
      POLYGON 1.645 0.305 1.645 0.115 1.43 0.115 1.43 0.165 1.595 0.165 1.595 0.305 ;
    LAYER M2 ;
      RECT 1.375 0.725 1.985 0.775 ;
    LAYER VIA1 ;
      RECT 1.805 0.725 1.935 0.775 ;
      RECT 1.425 0.725 1.475 0.775 ;
  END
END XOR3_X0P7M_A12TUL_C35

MACRO NAND2_X0P7B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P7B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02135 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02135 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.05375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P7B_A12TUL_C35

MACRO NAND2_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.425 0.28 0.425 0.28 0.495 0.445 0.495 0.445 0.605 0.28 0.605 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0336 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.875 0.635 0.595 0.58 0.595 0.58 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0336 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.11 0.575 0.975 0.77 0.975 0.77 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.375 0.715 0.375 0.715 0.925 0.235 0.925 0.235 1.11 0.305 1.11 0.305 0.975 0.505 0.975 0.505 1.11 ;
    END
    ANTENNADIFFAREA 0.067 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 1.04 0.37 1.04 0.37 1.165 0.17 1.165 0.17 0.99 0.1 0.99 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X1P4M_A12TUL_C35

MACRO NAND2B_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2B_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.71 0.23 0.495 0.365 0.495 0.365 0.425 0.145 0.425 0.145 0.495 0.175 0.495 0.175 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011375 ;
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.365 0.725 0.365 0.575 0.31 0.575 0.31 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0336 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.11 0.71 0.975 0.905 0.975 0.905 0.325 0.565 0.325 0.565 0.175 0.515 0.175 0.515 0.375 0.85 0.375 0.85 0.925 0.37 0.925 0.37 1.11 0.44 1.11 0.44 0.975 0.64 0.975 0.64 1.11 ;
    END
    ANTENNADIFFAREA 0.067 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.85 1.165 0.85 1.03 0.77 1.03 0.77 1.165 0.575 1.165 0.575 1.04 0.505 1.04 0.505 1.165 0.305 1.165 0.305 0.95 0.235 0.95 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.175 1.045 0.175 0.965 0.075 0.965 0.075 0.375 0.415 0.375 0.415 0.575 0.65 0.575 0.65 0.505 0.465 0.505 0.465 0.325 0.16 0.325 0.16 0.105 0.11 0.105 0.11 0.325 0.025 0.325 0.025 1.045 ;
  END
END NAND2B_X1P4M_A12TUL_C35

MACRO AOI22BB_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22BB_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.625 1.005 0.625 1.005 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.955 0.525 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0637 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.31 0.605 1.31 0.325 0.845 0.325 0.845 0.605 0.9 0.605 0.9 0.375 1.255 0.375 1.255 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0637 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.615 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02975 ;
  END B0N
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.705 0.235 0.705 0.235 0.525 0.165 0.525 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02975 ;
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.915 0.7 0.775 1.445 0.775 1.445 0.225 1.105 0.225 1.105 0.095 1.055 0.095 1.055 0.225 0.71 0.225 0.71 0.095 0.64 0.095 0.64 0.275 1.39 0.275 1.39 0.725 0.65 0.725 0.65 0.915 ;
    END
    ANTENNADIFFAREA 0.126 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.355 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.775 0.035 0.775 0.165 0.845 0.165 0.845 0.035 1.31 0.035 1.31 0.17 1.39 0.17 1.39 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.835 1.035 0.835 0.875 1.055 0.875 1.055 1.005 1.105 1.005 1.105 0.875 1.325 0.875 1.325 1.02 1.375 1.02 1.375 0.825 0.785 0.825 0.785 0.985 0.565 0.985 0.565 0.845 0.515 0.845 0.515 1.035 ;
      POLYGON 0.43 1.015 0.43 0.875 0.465 0.875 0.465 0.595 0.785 0.595 0.785 0.525 0.465 0.525 0.465 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.415 0.375 0.415 0.825 0.38 0.825 0.38 1.015 ;
  END
END AOI22BB_X2M_A12TUL_C35

MACRO NAND2_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.675 0.53 0.525 0.33 0.525 0.33 0.475 0.5 0.475 0.5 0.425 0.28 0.425 0.28 0.575 0.48 0.575 0.48 0.625 0.415 0.625 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0476 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0476 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.045 0.565 0.875 0.77 0.875 0.77 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.045 0.295 1.045 0.295 0.875 0.515 0.875 0.515 1.045 ;
    END
    ANTENNADIFFAREA 0.095 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.87 0.1 0.87 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND2_X2M_A12TUL_C35

MACRO BUF_X11M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X11M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.16 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.98 0.7 0.885 0.92 0.885 0.92 0.965 0.97 0.965 0.97 0.885 1.19 0.885 1.19 0.965 1.24 0.965 1.24 0.885 1.46 0.885 1.46 0.965 1.51 0.965 1.51 0.885 1.73 0.885 1.73 0.965 1.78 0.965 1.78 0.885 2 0.885 2 0.965 2.05 0.965 2.05 0.885 2.135 0.885 2.135 0.315 2.05 0.315 2.05 0.235 2 0.235 2 0.315 1.78 0.315 1.78 0.235 1.73 0.235 1.73 0.315 1.51 0.315 1.51 0.235 1.46 0.235 1.46 0.315 1.24 0.315 1.24 0.235 1.19 0.235 1.19 0.315 0.97 0.315 0.97 0.235 0.92 0.235 0.92 0.315 0.7 0.315 0.7 0.22 0.65 0.22 0.65 0.41 2.04 0.41 2.04 0.79 0.65 0.79 0.65 0.98 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
      LAYER M1 ;
        POLYGON 2.16 1.235 2.16 1.165 1.925 1.165 1.925 0.945 1.855 0.945 1.855 1.165 1.655 1.165 1.655 0.945 1.585 0.945 1.585 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.945 1.045 0.945 1.045 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.16 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.355 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.585 0.035 1.585 0.255 1.655 0.255 1.655 0.035 1.855 0.035 1.855 0.255 1.925 0.255 1.925 0.035 2.16 0.035 2.16 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 2.16 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1 0.43 0.875 0.565 0.875 0.565 0.725 0.635 0.725 0.635 0.565 1.92 0.565 1.92 0.605 1.99 0.605 1.99 0.515 0.585 0.515 0.585 0.675 0.515 0.675 0.515 0.825 0.085 0.825 0.085 0.375 0.43 0.375 0.43 0.185 0.38 0.185 0.38 0.325 0.16 0.325 0.16 0.2 0.11 0.2 0.11 0.325 0.035 0.325 0.035 0.875 0.11 0.875 0.11 1 0.16 1 0.16 0.875 0.38 0.875 0.38 1 ;
  END
END BUF_X11M_A12TUL_C35

MACRO BUFH_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02835 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.175 0.38 0.175 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.655 0.525 0.655 0.525 0.585 0.425 0.585 0.425 0.595 0.28 0.595 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X1P4M_A12TUL_C35

MACRO INV_X0P8M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P8M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.058125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P8M_A12TUL_C35

MACRO NAND2XB_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2XB_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.014525 ;
  END BN
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.775 0.665 0.625 0.465 0.625 0.465 0.575 0.645 0.575 0.645 0.525 0.415 0.525 0.415 0.675 0.615 0.675 0.615 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0476 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.875 0.905 0.875 0.905 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.85 0.375 0.85 0.825 0.38 0.825 0.38 1.045 0.43 1.045 0.43 0.875 0.65 0.875 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.095 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.87 0.235 0.87 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.305 0.305 0.035 0.775 0.035 0.775 0.27 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.095 0.16 0.89 0.085 0.89 0.085 0.425 0.31 0.425 0.31 0.595 0.36 0.595 0.36 0.475 0.715 0.475 0.715 0.69 0.765 0.69 0.765 0.425 0.36 0.425 0.36 0.375 0.16 0.375 0.16 0.145 0.11 0.145 0.11 0.375 0.035 0.375 0.035 0.94 0.11 0.94 0.11 1.095 ;
  END
END NAND2XB_X2M_A12TUL_C35

MACRO AO21B_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21B_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.575 0.235 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.165 0.375 0.165 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.019775 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.445 0.31 0.445 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.019775 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.525 0.6 0.525 0.6 0.475 0.77 0.475 0.77 0.425 0.55 0.425 0.55 0.575 0.75 0.575 0.75 0.625 0.685 0.625 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0427 ;
  END B0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.7 0.325 0.7 0.175 0.65 0.175 0.65 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.093 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.265 0.44 0.265 0.44 0.035 0.91 0.035 0.91 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.02 0.295 0.875 0.465 0.875 0.465 0.775 0.9 0.775 0.9 0.56 0.85 0.56 0.85 0.725 0.495 0.725 0.495 0.565 0.445 0.565 0.445 0.725 0.415 0.725 0.415 0.825 0.075 0.825 0.075 0.275 0.17 0.275 0.17 0.095 0.1 0.095 0.1 0.225 0.025 0.225 0.025 0.875 0.245 0.875 0.245 1.02 ;
  END
END AO21B_X1P4M_A12TUL_C35

MACRO INV_X0P8B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P8B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02205 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.15 0.23 0.15 0.23 0.23 0.31 0.23 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.04725 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.21 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P8B_A12TUL_C35

MACRO INV_X0P7B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P7B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.295 0.23 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01855 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.045 0.295 0.905 0.365 0.905 0.365 0.125 0.23 0.125 0.23 0.205 0.31 0.205 0.31 0.855 0.245 0.855 0.245 1.045 ;
    END
    ANTENNADIFFAREA 0.03975 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.855 0.1 0.855 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.18 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P7B_A12TUL_C35

MACRO INV_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P7M_A12TUL_C35

MACRO AO21_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO21_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.675 0.665 0.605 0.5 0.605 0.5 0.465 0.445 0.465 0.445 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.017325 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.065 0.835 0.925 0.905 0.925 0.905 0.295 0.835 0.295 0.835 0.15 0.785 0.15 0.785 0.345 0.85 0.345 0.85 0.875 0.785 0.875 0.785 1.065 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.305 0.17 0.035 0.505 0.035 0.505 0.195 0.575 0.195 0.575 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.015 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.015 ;
      POLYGON 0.565 0.98 0.565 0.825 0.77 0.825 0.77 0.425 0.63 0.425 0.63 0.325 0.43 0.325 0.43 0.12 0.38 0.12 0.38 0.375 0.58 0.375 0.58 0.475 0.715 0.475 0.715 0.775 0.515 0.775 0.515 0.98 ;
  END
END AO21_X0P7M_A12TUL_C35

MACRO INV_X0P6B_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P6B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.295 0.23 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015575 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.045 0.295 0.905 0.365 0.905 0.365 0.1 0.23 0.1 0.23 0.18 0.31 0.18 0.31 0.855 0.245 0.855 0.245 1.045 ;
    END
    ANTENNADIFFAREA 0.033375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.855 0.1 0.855 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.18 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P6B_A12TUL_C35

MACRO NOR2_X1B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X1B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.38 0.635 0.38 0.425 0.145 0.425 0.145 0.475 0.3 0.475 0.3 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02205 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02205 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.225 0.305 0.225 0.305 0.1 0.235 0.1 0.235 0.275 0.445 0.275 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.05025 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.18 0.17 0.035 0.365 0.035 0.365 0.175 0.445 0.175 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.18 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X1B_A12TUL_C35

MACRO OAI31_X2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OAI31_X2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.8 0.675 0.8 0.525 0.6 0.525 0.6 0.475 0.77 0.475 0.77 0.425 0.55 0.425 0.55 0.575 0.75 0.575 0.75 0.625 0.685 0.625 0.685 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.5 0.725 0.5 0.495 0.445 0.495 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.31 0.775 1.31 0.525 1.09 0.525 1.09 0.575 1.255 0.575 1.255 0.725 1.09 0.725 1.09 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0476 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.24 1.045 1.24 0.875 1.445 0.875 1.445 0.325 1.25 0.325 1.25 0.195 1.18 0.195 1.18 0.375 1.39 0.375 1.39 0.825 0.64 0.825 0.64 1.005 0.71 1.005 0.71 0.875 1.19 0.875 1.19 1.045 ;
    END
    ANTENNADIFFAREA 0.119 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 1.385 1.165 1.385 0.93 1.315 0.93 1.315 1.165 1.115 1.165 1.115 0.93 1.045 0.93 1.045 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.255 0.845 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.98 1.115 0.98 0.93 0.91 0.93 0.91 1.065 0.43 1.065 0.43 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1.115 ;
      POLYGON 1.105 0.375 1.105 0.135 1.315 0.135 1.315 0.27 1.385 0.27 1.385 0.085 1.055 0.085 1.055 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OAI31_X2M_A12TUL_C35

MACRO AOI22_X3M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22_X3M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.89 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.495 0.85 0.495 0.85 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.8 0.605 0.8 0.525 0.635 0.525 0.635 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.04 0.705 1.04 0.475 1.39 0.475 1.39 0.605 1.61 0.605 1.61 0.525 1.445 0.525 1.445 0.425 0.985 0.425 0.985 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.715 0.775 1.715 0.49 1.66 0.49 1.66 0.725 1.325 0.725 1.325 0.525 1.09 0.525 1.09 0.605 1.255 0.605 1.255 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09135 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.115 1.005 1.115 0.875 1.325 0.875 1.325 1 1.375 1 1.375 0.875 1.595 0.875 1.595 1 1.645 1 1.645 0.875 1.85 0.875 1.85 0.325 1.51 0.325 1.51 0.2 1.46 0.2 1.46 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 1.795 0.375 1.795 0.825 1.045 0.825 1.045 1.005 ;
    END
    ANTENNADIFFAREA 0.261 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
      LAYER M1 ;
        POLYGON 1.89 1.235 1.89 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.89 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.355 0.17 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 1.18 0.035 1.18 0.255 1.25 0.255 1.25 0.035 1.72 0.035 1.72 0.27 1.79 0.27 1.79 0.035 1.89 0.035 1.89 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.89 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.79 1.115 1.79 0.925 1.72 0.925 1.72 1.065 1.51 1.065 1.51 0.94 1.46 0.94 1.46 1.065 1.24 1.065 1.24 0.94 1.19 0.94 1.19 1.065 0.97 1.065 0.97 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.38 0.875 0.38 1 0.43 1 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.92 0.875 0.92 1.115 ;
  END
END AOI22_X3M_A12TUL_C35

MACRO NOR2_X1P4A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X1P4A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.425 0.28 0.425 0.28 0.495 0.445 0.495 0.445 0.605 0.28 0.605 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04235 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.495 0.58 0.495 0.58 0.725 0.23 0.725 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04235 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.13 0.515 0.13 0.515 0.325 0.295 0.325 0.295 0.13 0.245 0.13 0.245 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.085 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NOR2_X1P4A_A12TUL_C35

MACRO BUFH_X1P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.0775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.6 0.525 0.6 0.525 0.53 0.425 0.53 0.425 0.54 0.28 0.54 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X1P7M_A12TUL_C35

MACRO ADDF_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN ADDF_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.565 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.725 0.625 0.855 0.675 ;
        RECT 1.39 0.625 1.44 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 0.9 0.675 0.9 0.505 0.85 0.505 0.85 0.625 0.495 0.625 0.495 0.505 0.445 0.505 0.445 0.675 ;
        POLYGON 1.47 0.675 1.47 0.605 1.45 0.605 1.45 0.415 1.38 0.415 1.38 0.605 1.36 0.605 1.36 0.675 ;
        POLYGON 1.995 0.725 1.995 0.535 1.925 0.535 1.925 0.625 1.785 0.625 1.785 0.675 1.925 0.675 1.925 0.725 ;
      LAYER M2 ;
        RECT 0.675 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.1071 LAYER M2 ;
    ANTENNAGATEAREA 0.1071 LAYER M3 ;
    ANTENNAGATEAREA 0.1071 LAYER M4 ;
    ANTENNAGATEAREA 0.1071 LAYER M5 ;
    ANTENNAGATEAREA 0.1071 LAYER M6 ;
    ANTENNAGATEAREA 0.1071 LAYER M7 ;
    ANTENNAGATEAREA 0.1071 LAYER M8 ;
    ANTENNAGATEAREA 0.1071 LAYER AP ;
    ANTENNAMAXAREACAR 1.288889 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.605 0.525 0.655 0.575 ;
        RECT 1.53 0.525 1.58 0.575 ;
        RECT 2.065 0.525 2.115 0.575 ;
      LAYER M1 ;
        RECT 0.565 0.505 0.785 0.575 ;
        RECT 1.525 0.415 1.595 0.685 ;
        RECT 2.065 0.435 2.115 0.755 ;
      LAYER M2 ;
        RECT 0.555 0.525 2.165 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.1071 LAYER M2 ;
    ANTENNAGATEAREA 0.1071 LAYER M3 ;
    ANTENNAGATEAREA 0.1071 LAYER M4 ;
    ANTENNAGATEAREA 0.1071 LAYER M5 ;
    ANTENNAGATEAREA 0.1071 LAYER M6 ;
    ANTENNAGATEAREA 0.1071 LAYER M7 ;
    ANTENNAGATEAREA 0.1071 LAYER M8 ;
    ANTENNAGATEAREA 0.1071 LAYER AP ;
    ANTENNAMAXAREACAR 1.015873 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1587302 LAYER VIA1 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.985 0.425 1.035 0.475 ;
        RECT 1.25 0.425 1.3 0.475 ;
        RECT 1.825 0.425 1.955 0.475 ;
      LAYER M1 ;
        POLYGON 1.855 0.565 1.855 0.475 1.995 0.475 1.995 0.425 1.785 0.425 1.785 0.565 ;
        POLYGON 1.045 0.675 1.045 0.495 1.065 0.495 1.065 0.425 0.955 0.425 0.955 0.495 0.975 0.495 0.975 0.675 ;
        POLYGON 1.31 0.675 1.31 0.495 1.33 0.495 1.33 0.425 1.22 0.425 1.22 0.495 1.24 0.495 1.24 0.675 ;
      LAYER M2 ;
        RECT 0.935 0.425 2.005 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.0749 LAYER M2 ;
    ANTENNAGATEAREA 0.0749 LAYER M3 ;
    ANTENNAGATEAREA 0.0749 LAYER M4 ;
    ANTENNAGATEAREA 0.0749 LAYER M5 ;
    ANTENNAGATEAREA 0.0749 LAYER M6 ;
    ANTENNAGATEAREA 0.0749 LAYER M7 ;
    ANTENNAGATEAREA 0.0749 LAYER M8 ;
    ANTENNAGATEAREA 0.0749 LAYER AP ;
    ANTENNAMAXAREACAR 1.066667 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.825 0.095 0.825 0.095 0.375 0.295 0.375 0.295 0.165 0.245 0.165 0.245 0.325 0.04 0.325 0.04 0.875 0.245 0.875 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.32 1.015 2.32 0.875 2.525 0.875 2.525 0.325 2.32 0.325 2.32 0.165 2.27 0.165 2.27 0.375 2.47 0.375 2.47 0.825 2.27 0.825 2.27 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
      LAYER M1 ;
        POLYGON 2.565 1.235 2.565 1.165 2.465 1.165 2.465 0.93 2.395 0.93 2.395 1.165 2.195 1.165 2.195 0.945 2.125 0.945 2.125 1.165 1.52 1.165 1.52 0.945 1.45 0.945 1.45 1.165 1.25 1.165 1.25 0.865 1.18 0.865 1.18 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.565 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.375 0.44 0.035 0.64 0.035 0.64 0.305 0.71 0.305 0.71 0.035 1.18 0.035 1.18 0.27 1.25 0.27 1.25 0.035 1.45 0.035 1.45 0.255 1.52 0.255 1.52 0.035 2.125 0.035 2.125 0.255 2.195 0.255 2.195 0.035 2.395 0.035 2.395 0.27 2.465 0.27 2.465 0.035 2.565 0.035 2.565 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.275 0.17 0.275 0.17 0.035 0.37 0.035 0.37 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.565 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.105 1.055 1.105 0.865 1.055 0.865 1.055 1.005 0.835 1.005 0.835 0.825 0.515 0.825 0.515 1.015 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1.055 ;
      POLYGON 1.78 1.035 1.78 0.895 2.22 0.895 2.22 0.595 2.405 0.595 2.405 0.525 2.22 0.525 2.22 0.315 1.78 0.315 1.78 0.175 1.73 0.175 1.73 0.365 2.17 0.365 2.17 0.845 1.73 0.845 1.73 1.035 ;
      POLYGON 1.645 1.035 1.645 0.845 1.325 0.845 1.325 1.035 1.375 1.035 1.375 0.895 1.595 0.895 1.595 1.035 ;
      POLYGON 0.97 0.9 0.97 0.775 1.12 0.775 1.12 0.795 1.71 0.795 1.71 0.47 1.66 0.47 1.66 0.745 1.17 0.745 1.17 0.325 0.98 0.325 0.98 0.195 0.91 0.195 0.91 0.375 1.12 0.375 1.12 0.725 0.36 0.725 0.36 0.505 0.16 0.505 0.16 0.575 0.31 0.575 0.31 0.775 0.92 0.775 0.92 0.9 ;
      POLYGON 0.835 0.425 0.835 0.135 1.045 0.135 1.045 0.27 1.115 0.27 1.115 0.085 0.785 0.085 0.785 0.375 0.565 0.375 0.565 0.235 0.515 0.235 0.515 0.425 ;
      POLYGON 1.645 0.355 1.645 0.165 1.595 0.165 1.595 0.305 1.375 0.305 1.375 0.165 1.325 0.165 1.325 0.355 ;
  END
END ADDF_X1P4M_A12TUL_C35

MACRO AOI22BB_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI22BB_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.485 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.675 1.175 0.625 1.005 0.625 1.005 0.575 1.205 0.575 1.205 0.425 1.09 0.425 1.09 0.475 1.155 0.475 1.155 0.525 0.955 0.525 0.955 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0448 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.31 0.605 1.31 0.325 0.845 0.325 0.845 0.605 0.9 0.605 0.9 0.375 1.255 0.375 1.255 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0448 ;
  END A1
  PIN B0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END B0N
  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.705 0.235 0.705 0.235 0.525 0.165 0.525 0.165 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0224 ;
  END B1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.955 0.7 0.775 1.445 0.775 1.445 0.225 1.105 0.225 1.105 0.095 1.055 0.095 1.055 0.225 0.71 0.225 0.71 0.095 0.64 0.095 0.64 0.275 1.39 0.275 1.39 0.725 0.65 0.725 0.65 0.955 ;
    END
    ANTENNADIFFAREA 0.0885 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
      LAYER M1 ;
        POLYGON 1.485 1.235 1.485 1.165 1.25 1.165 1.25 0.945 1.18 0.945 1.18 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.485 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.32 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.775 0.035 0.775 0.165 0.845 0.165 0.845 0.035 1.31 0.035 1.31 0.17 1.39 0.17 1.39 0.035 1.485 0.035 1.485 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.32 ;
      LAYER M2 ;
        RECT 0 -0.065 1.485 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.835 1.075 0.835 0.875 1.055 0.875 1.055 1.005 1.105 1.005 1.105 0.875 1.325 0.875 1.325 1.02 1.375 1.02 1.375 0.825 0.785 0.825 0.785 1.025 0.565 1.025 0.565 0.885 0.515 0.885 0.515 1.075 ;
      POLYGON 0.43 1.015 0.43 0.875 0.465 0.875 0.465 0.595 0.785 0.595 0.785 0.525 0.465 0.525 0.465 0.325 0.295 0.325 0.295 0.145 0.245 0.145 0.245 0.375 0.415 0.375 0.415 0.825 0.38 0.825 0.38 1.015 ;
  END
END AOI22BB_X1P4M_A12TUL_C35

MACRO AND3_X1P4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND3_X1P4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.69 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.015 0.7 0.875 0.905 0.875 0.905 0.325 0.7 0.325 0.7 0.175 0.65 0.175 0.65 0.375 0.85 0.375 0.85 0.825 0.65 0.825 0.65 1.015 ;
    END
    ANTENNADIFFAREA 0.065 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.06 0.43 1.06 0.43 0.875 0.6 0.875 0.6 0.68 0.785 0.68 0.785 0.61 0.55 0.61 0.55 0.825 0.075 0.825 0.075 0.335 0.16 0.335 0.16 0.145 0.11 0.145 0.11 0.285 0.025 0.285 0.025 0.875 0.11 0.875 0.11 1.07 ;
  END
END AND3_X1P4M_A12TUL_C35

MACRO MXIT2_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN MXIT2_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.215 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.07 0.875 1.07 0.805 0.905 0.805 0.905 0.515 0.85 0.515 0.85 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03185 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.705 0.23 0.705 0.23 0.495 0.175 0.495 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03185 ;
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.455 0.525 0.505 0.575 ;
        RECT 0.99 0.525 1.04 0.575 ;
      LAYER M1 ;
        RECT 0.98 0.395 1.05 0.705 ;
        RECT 0.445 0.495 0.515 0.755 ;
      LAYER M2 ;
        RECT 0.405 0.525 1.09 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 LAYER M1 ;
    ANTENNAGATEAREA 0.03605 LAYER M2 ;
    ANTENNAGATEAREA 0.03605 LAYER M3 ;
    ANTENNAGATEAREA 0.03605 LAYER M4 ;
    ANTENNAGATEAREA 0.03605 LAYER M5 ;
    ANTENNAGATEAREA 0.03605 LAYER M6 ;
    ANTENNAGATEAREA 0.03605 LAYER M7 ;
    ANTENNAGATEAREA 0.03605 LAYER M8 ;
    ANTENNAGATEAREA 0.03605 LAYER AP ;
    ANTENNAMAXAREACAR 1.441861 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.166113 LAYER VIA1 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.395 0.475 0.395 0.475 0.445 0.58 0.445 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.06 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
      LAYER M1 ;
        POLYGON 1.215 1.235 1.215 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.17 1.165 0.17 0.925 0.1 0.925 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.215 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.305 0.17 0.035 0.91 0.035 0.91 0.16 0.98 0.16 0.98 0.035 1.215 0.035 1.215 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 1.215 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.115 1.105 1.115 0.975 1.175 0.975 1.175 0.225 1.115 0.225 1.115 0.09 1.045 0.09 1.045 0.225 0.85 0.225 0.85 0.085 0.53 0.085 0.53 0.295 0.345 0.295 0.345 0.5 0.295 0.5 0.295 0.57 0.395 0.57 0.395 0.345 0.58 0.345 0.58 0.135 0.8 0.135 0.8 0.275 1.125 0.275 1.125 0.925 1.045 0.925 1.045 1.105 ;
      POLYGON 0.845 1.105 0.845 0.925 0.745 0.925 0.745 0.395 0.865 0.395 0.865 0.345 0.745 0.345 0.745 0.255 0.635 0.255 0.635 0.335 0.695 0.335 0.695 0.925 0.505 0.925 0.505 1.105 0.575 1.105 0.575 0.975 0.775 0.975 0.775 1.105 ;
      POLYGON 0.295 1.015 0.295 0.825 0.09 0.825 0.09 0.425 0.295 0.425 0.295 0.245 0.46 0.245 0.46 0.195 0.245 0.195 0.245 0.375 0.04 0.375 0.04 0.875 0.245 0.875 0.245 1.015 ;
  END
END MXIT2_X1M_A12TUL_C35

MACRO AND3_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND3_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0203 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.105 0.71 1.005 0.77 1.005 0.77 0.395 0.7 0.395 0.7 0.255 0.65 0.255 0.65 0.445 0.715 0.445 0.715 0.925 0.64 0.925 0.64 1.105 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.95 0.235 0.95 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.06 0.43 1.06 0.43 0.875 0.63 0.875 0.63 0.505 0.58 0.505 0.58 0.825 0.075 0.825 0.075 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.025 0.305 0.025 0.875 0.11 0.875 0.11 1.07 ;
  END
END AND3_X1M_A12TUL_C35

MACRO MXIT2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN MXIT2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.605 0.365 0.325 0.145 0.325 0.145 0.395 0.31 0.395 0.31 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02345 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.91 0.665 0.91 0.495 0.935 0.495 0.935 0.425 0.82 0.425 0.82 0.495 0.84 0.495 0.84 0.665 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02345 ;
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.175 0.625 0.225 0.675 ;
        RECT 0.58 0.625 0.63 0.675 ;
      LAYER M1 ;
        POLYGON 0.665 0.675 0.665 0.605 0.64 0.605 0.64 0.42 0.57 0.42 0.57 0.605 0.545 0.605 0.545 0.675 ;
        RECT 0.165 0.465 0.235 0.755 ;
      LAYER M2 ;
        RECT 0.125 0.625 0.68 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0126 LAYER M1 ;
    ANTENNAGATEAREA 0.02975 LAYER M2 ;
    ANTENNAGATEAREA 0.02975 LAYER M3 ;
    ANTENNAGATEAREA 0.02975 LAYER M4 ;
    ANTENNAGATEAREA 0.02975 LAYER M5 ;
    ANTENNAGATEAREA 0.02975 LAYER M6 ;
    ANTENNAGATEAREA 0.02975 LAYER M7 ;
    ANTENNAGATEAREA 0.02975 LAYER M8 ;
    ANTENNAGATEAREA 0.02975 LAYER AP ;
    ANTENNAMAXAREACAR 1.611111 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1984127 LAYER VIA1 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.005 0.71 0.875 1.04 0.875 1.04 0.2 0.825 0.2 0.825 0.085 0.5 0.085 0.5 0.165 0.58 0.165 0.58 0.135 0.775 0.135 0.775 0.25 0.985 0.25 0.985 0.825 0.64 0.825 0.64 1.005 ;
    END
    ANTENNADIFFAREA 0.049 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.985 1.165 0.985 0.935 0.905 0.935 0.905 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.89 0.035 0.89 0.15 1 0.15 1 0.1 0.96 0.1 0.96 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.795 1.115 0.795 1.065 0.43 1.065 0.43 0.825 0.09 0.825 0.09 0.235 0.175 0.235 0.175 0.155 0.04 0.155 0.04 0.875 0.11 0.875 0.11 0.975 0.16 0.975 0.16 0.875 0.38 0.875 0.38 1.115 ;
      POLYGON 0.565 0.955 0.565 0.725 0.495 0.725 0.495 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.725 0.35 0.725 0.35 0.775 0.515 0.775 0.515 0.955 ;
      POLYGON 0.865 0.775 0.865 0.725 0.765 0.725 0.765 0.35 0.865 0.35 0.865 0.3 0.715 0.3 0.715 0.19 0.635 0.19 0.635 0.35 0.715 0.35 0.715 0.775 ;
  END
END MXIT2_X0P7M_A12TUL_C35

MACRO AND2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AND2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.565 0.17 0.565 0.17 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01225 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01225 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0.17 1.165 0.17 1.01 0.1 1.01 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.09 0.295 0.875 0.495 0.875 0.495 0.325 0.17 0.325 0.17 0.09 0.1 0.09 0.1 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.09 ;
  END
END AND2_X0P7M_A12TUL_C35

MACRO BUFH_X3P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X3P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.525 0.145 0.525 0.145 0.575 0.345 0.575 0.345 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.5 0.775 0.5 0.565 0.84 0.565 0.84 0.605 0.91 0.605 0.91 0.515 0.45 0.515 0.45 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUFH_X3P5M_A12TUL_C35

MACRO OA22_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA22_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.555 0.23 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.17 0.375 0.17 0.555 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.545 0.575 0.545 0.575 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.98 1.105 0.98 1.005 1.04 1.005 1.04 0.195 0.98 0.195 0.98 0.095 0.91 0.095 0.91 0.275 0.985 0.275 0.985 0.925 0.91 0.925 0.91 1.105 ;
    END
    ANTENNADIFFAREA 0.04875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.85 1.165 0.85 0.93 0.77 0.93 0.77 1.165 0.715 1.165 0.715 0.93 0.635 0.93 0.635 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.015 0.43 0.875 0.905 0.875 0.905 0.325 0.565 0.325 0.565 0.205 0.515 0.205 0.515 0.375 0.85 0.375 0.85 0.825 0.38 0.825 0.38 1.015 ;
      POLYGON 0.43 0.275 0.43 0.135 0.64 0.135 0.64 0.27 0.71 0.27 0.71 0.085 0.38 0.085 0.38 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OA22_X0P7M_A12TUL_C35

MACRO BUFH_X3M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUFH_X3M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.525 0.145 0.525 0.145 0.575 0.345 0.575 0.345 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.05565 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 0.905 0.875 0.905 0.325 0.835 0.325 0.835 0.2 0.785 0.2 0.785 0.325 0.565 0.325 0.565 0.185 0.515 0.185 0.515 0.375 0.85 0.375 0.85 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.355 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 0.17 0.27 0.17 0.035 0.37 0.035 0.37 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.9 0.295 0.775 0.495 0.775 0.495 0.565 0.705 0.565 0.705 0.605 0.775 0.605 0.775 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.375 0.295 0.375 0.295 0.185 0.245 0.185 0.245 0.325 0.025 0.325 0.025 0.775 0.245 0.775 0.245 0.9 ;
  END
END BUFH_X3M_A12TL_C35

MACRO INV_X3M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X3M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.575 0.315 0.575 0.315 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.635 0.875 0.635 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.58 0.375 0.58 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.161 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END INV_X3M_A12TL_C35

MACRO INV_X2M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X2M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.395 0.575 0.395 0.425 0.28 0.425 0.28 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0644 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X2M_A12TL_C35

MACRO BUFH_X1P7M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1P7M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.0775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.6 0.525 0.6 0.525 0.53 0.425 0.53 0.425 0.54 0.28 0.54 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X1P7M_A12TL_C35

MACRO BUF_X2P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X2P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.023275 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.77 0.875 0.77 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.133875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.9 0.235 0.9 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.955 0.16 0.83 0.33 0.83 0.33 0.67 0.63 0.67 0.63 0.56 0.58 0.56 0.58 0.62 0.28 0.62 0.28 0.78 0.09 0.78 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.83 0.11 0.83 0.11 0.955 ;
  END
END BUF_X2P5M_A12TUL_C35

MACRO AO21A1AI2_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.03875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 1.005 0.64 1.005 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END AO21A1AI2_X0P5M_A12TL_C35

MACRO CGENI_X1M_A12TL_C35
  CLASS CORE ;
  FOREIGN CGENI_X1M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.495 0.58 0.495 0.58 0.625 0.24 0.625 0.24 0.525 0.16 0.525 0.16 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.575 0.53 0.505 0.365 0.505 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.005 0.71 0.875 0.905 0.875 0.905 0.325 0.71 0.325 0.71 0.195 0.64 0.195 0.64 0.375 0.85 0.375 0.85 0.825 0.64 0.825 0.64 1.005 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END CON
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.845 1.115 0.845 0.93 0.775 0.93 0.775 1.065 0.565 1.065 0.565 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.115 ;
      POLYGON 0.565 0.375 0.565 0.135 0.775 0.135 0.775 0.27 0.845 0.27 0.845 0.085 0.515 0.085 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 ;
  END
END CGENI_X1M_A12TL_C35

MACRO BUF_X1P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X1P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.0775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.065 0.16 0.825 0.33 0.825 0.33 0.675 0.515 0.675 0.515 0.605 0.28 0.605 0.28 0.775 0.09 0.775 0.09 0.27 0.17 0.27 0.17 0.09 0.1 0.09 0.1 0.22 0.04 0.22 0.04 0.825 0.11 0.825 0.11 1.065 ;
  END
END BUF_X1P7M_A12TUL_C35

MACRO BUFH_X1M_A12TL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.395 0.395 0.395 0.395 0.325 0.175 0.325 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021175 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.305 1.165 0.305 0.83 0.235 0.83 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.995 0.16 0.755 0.36 0.755 0.36 0.505 0.31 0.505 0.31 0.705 0.09 0.705 0.09 0.275 0.17 0.275 0.17 0.095 0.1 0.095 0.1 0.225 0.04 0.225 0.04 0.755 0.11 0.755 0.11 0.995 ;
  END
END BUFH_X1M_A12TL_C35

MACRO BUF_X0P7B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X0P7B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.395 0.395 0.395 0.395 0.325 0.175 0.325 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013125 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.905 0.5 0.905 0.5 0.125 0.365 0.125 0.365 0.205 0.445 0.205 0.445 0.855 0.38 0.855 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.0405 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.305 1.165 0.305 0.845 0.235 0.845 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.195 0.305 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.195 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.055 0.16 0.775 0.36 0.775 0.36 0.56 0.31 0.56 0.31 0.725 0.09 0.725 0.09 0.165 0.175 0.165 0.175 0.085 0.04 0.085 0.04 0.775 0.11 0.775 0.11 1.055 ;
  END
END BUF_X0P7B_A12TUL_C35

MACRO AOI22_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN AOI22_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.975 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.445 0.225 0.445 0.085 0.365 0.085 0.365 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.515 0.825 0.515 0.975 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.21 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.635 0.035 0.635 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X0P5M_A12TL_C35

MACRO NAND4_X0P5A_A12TUH_C35
  CLASS CORE ;
  FOREIGN NAND4_X0P5A_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.495 0.435 0.495 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.595 0.31 0.595 0.31 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.175 0.475 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.115 0.575 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.235 0.925 0.235 1.115 0.305 1.115 0.305 0.975 0.505 0.975 0.505 1.115 ;
    END
    ANTENNADIFFAREA 0.03675 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 1.04 0.37 1.04 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND4_X0P5A_A12TUH_C35

MACRO OA21A1OI2_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.525 0.235 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.165 0.375 0.165 0.525 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.635 0.505 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.56 0.575 0.56 0.575 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.07 0.7 0.93 0.77 0.93 0.77 0.225 0.575 0.225 0.575 0.09 0.505 0.09 0.505 0.275 0.715 0.275 0.715 0.88 0.65 0.88 0.65 1.07 ;
    END
    ANTENNADIFFAREA 0.037625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.17 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 0.305 0.165 0.305 0.035 0.635 0.035 0.635 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.515 0.875 0.515 1.06 0.565 1.06 0.565 0.825 0.11 0.825 0.11 1.07 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END OA21A1OI2_X0P5M_A12TL_C35

MACRO NAND2_X0P5A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P5A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.495 0.31 0.495 0.31 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.175 0.375 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.075 0.295 0.975 0.5 0.975 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.925 0.245 0.925 0.245 1.075 ;
    END
    ANTENNADIFFAREA 0.03125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.445 1.165 0.445 1.03 0.365 1.03 0.365 1.165 0.17 1.165 0.17 0.995 0.1 0.995 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P5A_A12TUL_C35

MACRO BUFH_X1P2M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X1P2M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02485 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.13 0.38 0.13 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.055 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.27 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.985 0.16 0.855 0.33 0.855 0.33 0.705 0.495 0.705 0.495 0.515 0.445 0.515 0.445 0.655 0.28 0.655 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.985 ;
  END
END BUFH_X1P2M_A12TUL_C35

MACRO NAND2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.495 0.31 0.495 0.31 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.175 0.375 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.04 0.295 0.975 0.5 0.975 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.925 0.245 0.925 0.245 1.04 ;
    END
    ANTENNADIFFAREA 0.04075 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.445 1.165 0.445 1.03 0.365 1.03 0.365 1.165 0.17 1.165 0.17 0.99 0.1 0.99 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P7M_A12TUL_C35

MACRO INV_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN INV_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.065 0.295 0.925 0.365 0.925 0.365 0.195 0.305 0.195 0.305 0.09 0.235 0.09 0.235 0.27 0.31 0.27 0.31 0.875 0.245 0.875 0.245 1.065 ;
    END
    ANTENNADIFFAREA 0.03525 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P5M_A12TUL_C35

MACRO OAI21_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN OAI21_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.565 0.3 0.565 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.635 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01295 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.065 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.065 ;
    END
    ANTENNADIFFAREA 0.03925 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 1 0.505 1 0.505 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END OAI21_X0P5M_A12TL_C35

MACRO AOI22_X0P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN AOI22_X0P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.975 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.445 0.225 0.445 0.085 0.365 0.085 0.365 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.515 0.825 0.515 0.975 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.21 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.635 0.035 0.635 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X0P5M_A12TH_C35

MACRO MXIT2_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN MXIT2_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.495 0.31 0.495 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.705 0.77 0.495 0.8 0.495 0.8 0.425 0.685 0.425 0.685 0.495 0.71 0.495 0.71 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02065 ;
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.55 0.63 0.55 0.63 0.44 0.58 0.44 0.58 0.495 0.445 0.495 0.445 0.725 0.23 0.725 0.23 0.565 0.175 0.565 0.175 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03395 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 0.975 0.715 0.975 0.715 0.875 0.905 0.875 0.905 0.325 0.71 0.325 0.71 0.225 0.575 0.225 0.575 0.095 0.505 0.095 0.505 0.275 0.66 0.275 0.66 0.375 0.85 0.375 0.85 0.825 0.665 0.825 0.665 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.059 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.845 1.165 0.845 0.93 0.775 0.93 0.775 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.845 0.27 0.845 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.775 0.035 0.775 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.05 0.16 0.875 0.61 0.875 0.61 0.735 0.65 0.735 0.65 0.665 0.56 0.665 0.56 0.825 0.085 0.825 0.085 0.375 0.445 0.375 0.445 0.435 0.495 0.435 0.495 0.325 0.16 0.325 0.16 0.15 0.11 0.15 0.11 0.325 0.035 0.325 0.035 0.875 0.11 0.875 0.11 1.05 ;
  END
END MXIT2_X0P5M_A12TL_C35

MACRO BUFH_X5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.35 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.195 0.625 0.195 0.575 0.53 0.575 0.53 0.425 0.415 0.425 0.415 0.475 0.48 0.475 0.48 0.525 0.145 0.525 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.092925 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.015 0.7 0.875 0.92 0.875 0.92 1 0.97 1 0.97 0.875 1.19 0.875 1.19 1 1.24 1 1.24 0.875 1.31 0.875 1.31 0.325 1.24 0.325 1.24 0.2 1.19 0.2 1.19 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.7 0.325 0.7 0.185 0.65 0.185 0.65 0.375 1.255 0.375 1.255 0.825 0.65 0.825 0.65 1.015 ;
    END
    ANTENNADIFFAREA 0.253 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
      LAYER M1 ;
        POLYGON 1.35 1.235 1.35 1.165 1.115 1.165 1.115 0.945 1.045 0.945 1.045 1.165 0.845 1.165 0.845 0.945 0.775 0.945 0.775 1.165 0.575 1.165 0.575 0.845 0.505 0.845 0.505 1.165 0.305 1.165 0.305 0.845 0.235 0.845 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.35 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.355 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.35 0.035 1.35 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 1.35 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.9 0.43 0.775 0.63 0.775 0.63 0.565 1.11 0.565 1.11 0.605 1.18 0.605 1.18 0.515 0.58 0.515 0.58 0.725 0.085 0.725 0.085 0.375 0.43 0.375 0.43 0.185 0.38 0.185 0.38 0.325 0.16 0.325 0.16 0.2 0.11 0.2 0.11 0.325 0.035 0.325 0.035 0.775 0.11 0.775 0.11 0.9 0.16 0.9 0.16 0.775 0.38 0.775 0.38 0.9 ;
  END
END BUFH_X5M_A12TUL_C35

MACRO INV_X4M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X4M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.675 0.5 0.575 0.665 0.575 0.665 0.425 0.55 0.425 0.55 0.475 0.615 0.475 0.615 0.525 0.145 0.525 0.145 0.575 0.45 0.575 0.45 0.625 0.28 0.625 0.28 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1 0.565 1 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.2 0.515 0.2 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 0.715 0.375 0.715 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.93 0.64 0.93 0.64 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.64 0.035 0.64 0.27 0.71 0.27 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END INV_X4M_A12TL_C35

MACRO NOR2_X0P5A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.295 0.225 0.295 0.145 0.245 0.145 0.245 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.205 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.205 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5A_A12TUL_C35

MACRO NAND2_X1B_A12TL_C35
  CLASS CORE ;
  FOREIGN NAND2_X1B_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0301 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.095 0.37 0.095 0.37 0.275 0.445 0.275 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.07575 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X1B_A12TL_C35

MACRO NOR2_X0P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.54 0.175 0.54 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0168 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.31 0.225 0.31 0.085 0.23 0.085 0.23 0.165 0.26 0.165 0.26 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.0385 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 0.17 0.17 0.17 0.035 0.365 0.035 0.365 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5B_A12TUL_C35

MACRO NOR2_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.31 0.225 0.31 0.095 0.23 0.095 0.23 0.175 0.26 0.175 0.26 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.030125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.175 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.175 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5M_A12TUH_C35

MACRO NAND2_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.495 0.31 0.495 0.31 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01225 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.605 0.23 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.175 0.375 0.175 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01225 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.09 0.295 0.975 0.5 0.975 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.925 0.245 0.925 0.245 1.09 ;
    END
    ANTENNADIFFAREA 0.02975 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.445 1.165 0.445 1.03 0.365 1.03 0.365 1.165 0.17 1.165 0.17 1.01 0.1 1.01 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P5M_A12TUL_C35

MACRO INV_X0P6M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X0P6M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01925 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.065 0.295 0.925 0.365 0.925 0.365 0.26 0.295 0.26 0.295 0.12 0.245 0.12 0.245 0.31 0.31 0.31 0.31 0.875 0.245 0.875 0.245 1.065 ;
    END
    ANTENNADIFFAREA 0.04125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.875 0.1 0.875 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.3 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.3 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P6M_A12TL_C35

MACRO ADDF_X1M_A12TL_C35
  CLASS CORE ;
  FOREIGN ADDF_X1M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.295 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.595 0.625 0.725 0.675 ;
        RECT 1.255 0.625 1.305 0.675 ;
        RECT 1.825 0.625 1.955 0.675 ;
      LAYER M1 ;
        POLYGON 0.765 0.675 0.765 0.505 0.715 0.505 0.715 0.625 0.36 0.625 0.36 0.505 0.31 0.505 0.31 0.675 ;
        POLYGON 1.335 0.675 1.335 0.605 1.315 0.605 1.315 0.415 1.245 0.415 1.245 0.605 1.225 0.605 1.225 0.675 ;
        POLYGON 1.855 0.725 1.855 0.675 2 0.675 2 0.625 1.855 0.625 1.855 0.535 1.785 0.535 1.785 0.725 ;
      LAYER M2 ;
        RECT 0.545 0.625 2.005 0.675 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.10465 LAYER M2 ;
    ANTENNAGATEAREA 0.10465 LAYER M3 ;
    ANTENNAGATEAREA 0.10465 LAYER M4 ;
    ANTENNAGATEAREA 0.10465 LAYER M5 ;
    ANTENNAGATEAREA 0.10465 LAYER M6 ;
    ANTENNAGATEAREA 0.10465 LAYER M7 ;
    ANTENNAGATEAREA 0.10465 LAYER M8 ;
    ANTENNAGATEAREA 0.10465 LAYER AP ;
    ANTENNAMAXAREACAR 1.304762 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.475 0.425 0.605 0.475 ;
        RECT 1.425 0.425 1.555 0.475 ;
        RECT 1.825 0.425 1.955 0.475 ;
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.425 0.435 0.425 0.435 0.575 0.505 0.575 0.505 0.475 0.575 0.475 0.575 0.575 ;
        POLYGON 1.995 0.575 1.995 0.425 1.785 0.425 1.785 0.475 1.925 0.475 1.925 0.575 ;
        POLYGON 1.455 0.605 1.455 0.475 1.595 0.475 1.595 0.425 1.385 0.425 1.385 0.605 ;
      LAYER M2 ;
        RECT 0.425 0.425 2.005 0.475 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.10465 LAYER M2 ;
    ANTENNAGATEAREA 0.10465 LAYER M3 ;
    ANTENNAGATEAREA 0.10465 LAYER M4 ;
    ANTENNAGATEAREA 0.10465 LAYER M5 ;
    ANTENNAGATEAREA 0.10465 LAYER M6 ;
    ANTENNAGATEAREA 0.10465 LAYER M7 ;
    ANTENNAGATEAREA 0.10465 LAYER M8 ;
    ANTENNAGATEAREA 0.10465 LAYER AP ;
    ANTENNAMAXAREACAR 1.111111 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.4126985 LAYER VIA1 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.85 0.525 0.9 0.575 ;
        RECT 1.11 0.525 1.16 0.575 ;
        RECT 1.665 0.525 1.715 0.575 ;
      LAYER M1 ;
        RECT 0.84 0.42 0.91 0.675 ;
        RECT 1.1 0.415 1.17 0.685 ;
        RECT 1.665 0.445 1.715 0.755 ;
      LAYER M2 ;
        RECT 0.8 0.525 1.765 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01575 LAYER M1 ;
    ANTENNAGATEAREA 0.07245 LAYER M2 ;
    ANTENNAGATEAREA 0.07245 LAYER M3 ;
    ANTENNAGATEAREA 0.07245 LAYER M4 ;
    ANTENNAGATEAREA 0.07245 LAYER M5 ;
    ANTENNAGATEAREA 0.07245 LAYER M6 ;
    ANTENNAGATEAREA 0.07245 LAYER M7 ;
    ANTENNAGATEAREA 0.07245 LAYER M8 ;
    ANTENNAGATEAREA 0.07245 LAYER AP ;
    ANTENNAMAXAREACAR 0.984127 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1587302 LAYER VIA1 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.17 1.105 0.17 0.925 0.095 0.925 0.095 0.27 0.17 0.27 0.17 0.09 0.1 0.09 0.1 0.195 0.04 0.195 0.04 1.005 0.1 1.005 0.1 1.105 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.195 1.105 2.195 1.005 2.255 1.005 2.255 0.195 2.195 0.195 2.195 0.09 2.125 0.09 2.125 0.27 2.2 0.27 2.2 0.925 2.125 0.925 2.125 1.105 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
      LAYER M1 ;
        POLYGON 2.295 1.235 2.295 1.165 2.06 1.165 2.06 0.905 1.99 0.905 1.99 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 1.115 1.165 1.115 0.855 1.045 0.855 1.045 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.855 0.235 0.855 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.295 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.375 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 1.045 0.035 1.045 0.27 1.115 0.27 1.115 0.035 1.315 0.035 1.315 0.255 1.385 0.255 1.385 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.295 0.035 2.295 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.375 ;
      LAYER M2 ;
        RECT 0 -0.065 2.295 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.97 1.065 0.97 0.875 0.92 0.875 0.92 1.015 0.7 1.015 0.7 0.845 0.38 0.845 0.38 1.035 0.43 1.035 0.43 0.895 0.65 0.895 0.65 1.065 ;
      POLYGON 1.645 1.045 1.645 0.905 1.845 0.905 1.845 0.835 2.12 0.835 2.12 0.325 1.645 0.325 1.645 0.165 1.595 0.165 1.595 0.375 2.07 0.375 2.07 0.785 1.795 0.785 1.795 0.855 1.595 0.855 1.595 1.045 ;
      POLYGON 1.51 1.035 1.51 0.845 1.19 0.845 1.19 1.035 1.24 1.035 1.24 0.895 1.46 0.895 1.46 1.035 ;
      POLYGON 0.835 0.91 0.835 0.785 1.58 0.785 1.58 0.605 1.53 0.605 1.53 0.735 1.035 0.735 1.035 0.32 0.845 0.32 0.845 0.19 0.775 0.19 0.775 0.37 0.985 0.37 0.985 0.735 0.225 0.735 0.225 0.505 0.175 0.505 0.175 0.785 0.785 0.785 0.785 0.91 ;
      POLYGON 0.7 0.375 0.7 0.135 0.91 0.135 0.91 0.27 0.98 0.27 0.98 0.085 0.65 0.085 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 ;
      POLYGON 1.51 0.355 1.51 0.165 1.46 0.165 1.46 0.305 1.24 0.305 1.24 0.165 1.19 0.165 1.19 0.355 ;
  END
END ADDF_X1M_A12TL_C35

MACRO AO1B2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AO1B2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.675 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011725 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.525 0.3 0.525 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011725 ;
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02135 ;
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 0.975 0.77 0.975 0.77 0.295 0.7 0.295 0.7 0.155 0.65 0.155 0.65 0.345 0.715 0.345 0.715 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.05375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 0.935 0.37 0.935 0.37 1.165 0.17 1.165 0.17 0.995 0.1 0.995 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.31 1.115 0.31 0.875 0.63 0.875 0.63 0.6 0.58 0.6 0.58 0.825 0.075 0.825 0.075 0.2 0.19 0.2 0.19 0.15 0.025 0.15 0.025 0.875 0.23 0.875 0.23 1.115 ;
  END
END AO1B2_X0P7M_A12TUL_C35

MACRO NOR2_X0P7B_A12TUL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P7B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.635 0.375 0.425 0.145 0.425 0.145 0.475 0.305 0.475 0.305 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018375 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.785 0.365 0.735 0.24 0.735 0.24 0.535 0.16 0.535 0.16 0.735 0.145 0.735 0.145 0.785 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018375 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.31 0.225 0.31 0.085 0.23 0.085 0.23 0.165 0.26 0.165 0.26 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.041875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.17 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P7B_A12TUL_C35

MACRO INV_X1M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X1M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.055 0.295 0.915 0.365 0.915 0.365 0.285 0.295 0.285 0.295 0.145 0.245 0.145 0.245 0.335 0.31 0.335 0.31 0.865 0.245 0.865 0.245 1.055 ;
    END
    ANTENNADIFFAREA 0.069 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.865 0.1 0.865 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X1M_A12TL_C35

MACRO NAND2_X0P5B_A12TL_C35
  CLASS CORE ;
  FOREIGN NAND2_X0P5B_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.695 0.365 0.495 0.31 0.495 0.31 0.625 0.145 0.625 0.145 0.695 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.09 0.295 0.875 0.5 0.875 0.5 0.195 0.44 0.195 0.44 0.09 0.37 0.09 0.37 0.27 0.445 0.27 0.445 0.825 0.245 0.825 0.245 1.09 ;
    END
    ANTENNADIFFAREA 0.03825 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.915 0.1 0.915 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NAND2_X0P5B_A12TL_C35

MACRO AOI211_X0P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN AOI211_X0P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021525 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.045 0.7 0.905 0.77 0.905 0.77 0.225 0.715 0.225 0.715 0.085 0.635 0.085 0.635 0.225 0.44 0.225 0.44 0.095 0.37 0.095 0.37 0.275 0.715 0.275 0.715 0.855 0.65 0.855 0.65 1.045 ;
    END
    ANTENNADIFFAREA 0.056125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.335 0.17 0.035 0.505 0.035 0.505 0.165 0.575 0.165 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.335 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 1.02 0.43 0.825 0.11 0.825 0.11 1.02 0.16 1.02 0.16 0.875 0.38 0.875 0.38 1.02 ;
  END
END AOI211_X0P5M_A12TUL_C35

MACRO BUF_X4B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X4B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.04 0.875 1.04 0.325 0.835 0.325 0.835 0.095 0.785 0.095 0.785 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.375 0.985 0.375 0.985 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.144 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.31 0.305 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.27 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.31 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 1.02 0.295 0.775 0.495 0.775 0.495 0.565 0.84 0.565 0.84 0.605 0.91 0.605 0.91 0.515 0.445 0.515 0.445 0.725 0.075 0.725 0.075 0.315 0.16 0.315 0.16 0.115 0.11 0.115 0.11 0.265 0.025 0.265 0.025 0.775 0.245 0.775 0.245 1.02 ;
  END
END BUF_X4B_A12TUL_C35

MACRO DLYCLK8S2_X2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN DLYCLK8S2_X2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 3.375 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.595 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0483 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 3.13 0.915 3.13 0.775 3.335 0.775 3.335 0.325 3.13 0.325 3.13 0.145 3.08 0.145 3.08 0.375 3.28 0.375 3.28 0.725 3.08 0.725 3.08 0.915 ;
    END
    ANTENNADIFFAREA 0.078 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
        RECT 2.405 1.175 2.455 1.225 ;
        RECT 2.54 1.175 2.59 1.225 ;
        RECT 2.675 1.175 2.725 1.225 ;
        RECT 2.81 1.175 2.86 1.225 ;
        RECT 2.945 1.175 2.995 1.225 ;
        RECT 3.08 1.175 3.13 1.225 ;
        RECT 3.215 1.175 3.265 1.225 ;
      LAYER M1 ;
        POLYGON 3.375 1.235 3.375 1.165 3.275 1.165 3.275 0.845 3.205 0.845 3.205 1.165 3.005 1.165 3.005 0.845 2.935 0.845 2.935 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 3.375 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
        RECT 2.405 -0.025 2.455 0.025 ;
        RECT 2.54 -0.025 2.59 0.025 ;
        RECT 2.675 -0.025 2.725 0.025 ;
        RECT 2.81 -0.025 2.86 0.025 ;
        RECT 2.945 -0.025 2.995 0.025 ;
        RECT 3.08 -0.025 3.13 0.025 ;
        RECT 3.215 -0.025 3.265 0.025 ;
      LAYER M1 ;
        POLYGON 3.275 0.27 3.275 0.035 3.375 0.035 3.375 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.37 0.035 0.37 0.21 0.44 0.21 0.44 0.035 2.935 0.035 2.935 0.27 3.005 0.27 3.005 0.035 3.205 0.035 3.205 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 3.375 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.73 0.575 2.8 1.065 ;
      RECT 2.595 0.575 2.665 1.065 ;
      RECT 2.46 0.575 2.53 1.065 ;
      RECT 2.325 0.575 2.395 1.065 ;
      RECT 2.19 0.575 2.26 1.065 ;
      RECT 2.055 0.575 2.125 1.065 ;
      RECT 1.92 0.575 1.99 1.065 ;
      RECT 1.785 0.575 1.855 1.065 ;
      RECT 1.65 0.575 1.72 1.065 ;
      RECT 1.515 0.575 1.585 1.065 ;
      RECT 1.38 0.575 1.45 1.065 ;
      RECT 1.245 0.575 1.315 1.065 ;
      RECT 1.11 0.575 1.18 1.065 ;
      RECT 0.975 0.575 1.045 1.065 ;
      RECT 0.84 0.575 0.91 1.065 ;
      RECT 0.705 0.575 0.775 1.065 ;
      RECT 0.57 0.575 0.64 1.065 ;
      POLYGON 0.295 0.915 0.295 0.775 0.495 0.775 0.495 0.475 2.995 0.475 2.995 0.585 3.075 0.585 3.075 0.475 3.135 0.475 3.135 0.585 3.215 0.585 3.215 0.425 0.495 0.425 0.495 0.28 0.31 0.28 0.31 0.095 0.23 0.095 0.23 0.33 0.445 0.33 0.445 0.725 0.245 0.725 0.245 0.915 ;
      POLYGON 2.8 0.325 2.8 0.135 2.73 0.135 2.73 0.275 2.665 0.275 2.665 0.135 2.595 0.135 2.595 0.275 2.53 0.275 2.53 0.135 2.46 0.135 2.46 0.275 2.395 0.275 2.395 0.135 2.325 0.135 2.325 0.275 2.26 0.275 2.26 0.135 2.19 0.135 2.19 0.275 2.125 0.275 2.125 0.135 2.055 0.135 2.055 0.275 1.99 0.275 1.99 0.135 1.92 0.135 1.92 0.275 1.855 0.275 1.855 0.135 1.785 0.135 1.785 0.275 1.72 0.275 1.72 0.135 1.65 0.135 1.65 0.275 1.585 0.275 1.585 0.135 1.515 0.135 1.515 0.275 1.45 0.275 1.45 0.135 1.38 0.135 1.38 0.275 1.315 0.275 1.315 0.135 1.245 0.135 1.245 0.275 1.18 0.275 1.18 0.135 1.11 0.135 1.11 0.275 1.045 0.275 1.045 0.135 0.975 0.135 0.975 0.275 0.91 0.275 0.91 0.135 0.84 0.135 0.84 0.275 0.775 0.275 0.775 0.135 0.705 0.135 0.705 0.275 0.64 0.275 0.64 0.135 0.57 0.135 0.57 0.325 ;
  END
END DLYCLK8S2_X2B_A12TUL_C35

MACRO INV_X1P2M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X1P2M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0385 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.015 0.295 0.875 0.5 0.875 0.5 0.325 0.295 0.325 0.295 0.13 0.245 0.13 0.245 0.375 0.445 0.375 0.445 0.825 0.245 0.825 0.245 1.015 ;
    END
    ANTENNADIFFAREA 0.055 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.44 1.165 0.44 0.93 0.37 0.93 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.305 0.17 0.035 0.37 0.035 0.37 0.27 0.44 0.27 0.44 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.305 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END INV_X1P2M_A12TL_C35

MACRO AOI21_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN AOI21_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.575 0.37 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.3 0.375 0.3 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.425 0.165 0.425 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.775 0.5 0.495 0.445 0.495 0.445 0.725 0.28 0.725 0.28 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.905 0.635 0.905 0.635 0.225 0.43 0.225 0.43 0.14 0.38 0.14 0.38 0.275 0.58 0.275 0.58 0.855 0.515 0.855 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.035375 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.21 0.17 0.035 0.5 0.035 0.5 0.17 0.58 0.17 0.58 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.065 0.43 1.065 0.43 0.825 0.11 0.825 0.11 1.07 ;
  END
END AOI21_X0P5M_A12TL_C35

MACRO OAI21_X0P7M_A12TL_C35
  CLASS CORE ;
  FOREIGN OAI21_X0P7M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.37 0.725 0.37 0.565 0.3 0.565 0.3 0.725 0.15 0.725 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.635 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.605 0.5 0.325 0.28 0.325 0.28 0.375 0.445 0.375 0.445 0.605 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01785 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.095 0.505 0.095 0.505 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.05425 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.58 1.165 0.58 0.93 0.5 0.93 0.5 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.095 0.37 0.095 0.37 0.225 0.17 0.225 0.17 0.095 0.1 0.095 0.1 0.275 ;
  END
END OAI21_X0P7M_A12TL_C35

MACRO NAND4BB_X0P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN NAND4BB_X0P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.725 0.235 0.575 0.365 0.575 0.365 0.525 0.145 0.525 0.145 0.575 0.165 0.575 0.165 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.665 0.31 0.665 0.31 0.805 0.15 0.805 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.675 0.645 0.425 0.415 0.425 0.415 0.475 0.565 0.475 0.565 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.565 0.435 0.565 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.095 0.835 0.975 0.905 0.975 0.905 0.195 0.845 0.195 0.845 0.09 0.775 0.09 0.775 0.27 0.85 0.27 0.85 0.925 0.515 0.925 0.515 1.085 0.565 1.085 0.565 0.975 0.785 0.975 0.785 1.095 ;
    END
    ANTENNADIFFAREA 0.041125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 1.035 0.64 1.035 0.64 1.165 0.44 1.165 0.44 0.94 0.37 0.94 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.11 0.17 0.93 0.075 0.93 0.075 0.375 0.715 0.375 0.715 0.515 0.77 0.515 0.77 0.325 0.305 0.325 0.305 0.09 0.235 0.09 0.235 0.325 0.025 0.325 0.025 0.98 0.1 0.98 0.1 1.11 ;
  END
END NAND4BB_X0P5M_A12TH_C35

MACRO NOR2_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.31 0.225 0.31 0.095 0.23 0.095 0.23 0.175 0.26 0.175 0.26 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.030125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.175 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.175 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5M_A12TL_C35

MACRO NOR4BB_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN NOR4BB_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0084 ;
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.395 0.31 0.395 0.31 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0084 ;
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.775 0.64 0.565 0.57 0.565 0.57 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.635 0.505 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.435 0.495 0.435 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.845 1.105 0.845 1.005 0.905 1.005 0.905 0.225 0.85 0.225 0.85 0.085 0.77 0.085 0.77 0.225 0.575 0.225 0.575 0.09 0.505 0.09 0.505 0.275 0.85 0.275 0.85 0.925 0.775 0.925 0.775 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.185 0.44 0.035 0.64 0.035 0.64 0.165 0.71 0.165 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.185 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.31 1.105 0.31 1.025 0.28 1.025 0.28 0.875 0.765 0.875 0.765 0.665 0.715 0.665 0.715 0.825 0.085 0.825 0.085 0.175 0.19 0.175 0.19 0.125 0.035 0.125 0.035 0.875 0.23 0.875 0.23 1.105 ;
  END
END NOR4BB_X0P5M_A12TUH_C35

MACRO AOI22_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN AOI22_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.55 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.31 0.375 0.31 0.55 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.975 0.565 0.875 0.77 0.875 0.77 0.325 0.565 0.325 0.565 0.225 0.445 0.225 0.445 0.085 0.365 0.085 0.365 0.275 0.515 0.275 0.515 0.375 0.715 0.375 0.715 0.825 0.515 0.825 0.515 0.975 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.715 0.21 0.715 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.21 0.17 0.21 0.17 0.035 0.635 0.035 0.635 0.21 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.71 1.11 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.11 ;
  END
END AOI22_X0P5M_A12TUH_C35

MACRO NAND3_X0P7A_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND3_X0P7A_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.705 0.5 0.425 0.28 0.425 0.28 0.475 0.445 0.475 0.445 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0175 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.37 0.825 0.37 0.625 0.3 0.625 0.3 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0175 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.775 0.235 0.575 0.365 0.575 0.365 0.525 0.145 0.525 0.145 0.575 0.165 0.575 0.165 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0175 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.11 0.575 0.975 0.635 0.975 0.635 0.295 0.565 0.295 0.565 0.155 0.515 0.155 0.515 0.345 0.58 0.345 0.58 0.925 0.235 0.925 0.235 1.11 0.305 1.11 0.305 0.975 0.505 0.975 0.505 1.11 ;
    END
    ANTENNADIFFAREA 0.0585 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.44 1.165 0.44 1.035 0.37 1.035 0.37 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.35 0.17 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.35 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END NAND3_X0P7A_A12TUL_C35

MACRO BUF_X2B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X2B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.325 0.43 0.325 0.43 0.095 0.38 0.095 0.38 0.375 0.58 0.375 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.072 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.27 0.575 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.27 0.305 0.27 0.305 0.035 0.505 0.035 0.505 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.995 0.16 0.825 0.33 0.825 0.33 0.595 0.515 0.595 0.515 0.525 0.425 0.525 0.425 0.535 0.28 0.535 0.28 0.775 0.09 0.775 0.09 0.19 0.175 0.19 0.175 0.11 0.04 0.11 0.04 0.825 0.11 0.825 0.11 0.995 ;
  END
END BUF_X2B_A12TUL_C35

MACRO AND4_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN AND4_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.625 0.235 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.165 0.475 0.165 0.625 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.775 0.395 0.725 0.365 0.725 0.365 0.595 0.31 0.595 0.31 0.705 0.15 0.705 0.15 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.505 0.625 0.505 0.495 0.435 0.495 0.435 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.07 0.835 0.93 0.905 0.93 0.905 0.195 0.845 0.195 0.845 0.085 0.775 0.085 0.775 0.27 0.85 0.27 0.85 0.88 0.785 0.88 0.785 1.07 ;
    END
    ANTENNADIFFAREA 0.034875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 0.885 0.64 0.885 0.64 1.165 0.44 1.165 0.44 1.005 0.37 1.005 0.37 1.165 0.17 1.165 0.17 1.005 0.1 1.005 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.71 0.255 0.71 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.64 0.035 0.64 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.08 0.565 0.815 0.765 0.815 0.765 0.625 0.715 0.625 0.715 0.765 0.515 0.765 0.515 0.86 0.085 0.86 0.085 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.035 0.305 0.035 0.91 0.245 0.91 0.245 1.08 0.295 1.08 0.295 0.91 0.515 0.91 0.515 1.08 ;
  END
END AND4_X0P5M_A12TUH_C35

MACRO BUF_X2P5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X2P5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018725 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.77 0.875 0.77 0.325 0.7 0.325 0.7 0.135 0.65 0.135 0.65 0.325 0.43 0.325 0.43 0.145 0.38 0.145 0.38 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.205 0.305 0.205 0.305 0.035 0.505 0.035 0.505 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.95 0.16 0.825 0.33 0.825 0.33 0.67 0.63 0.67 0.63 0.56 0.58 0.56 0.58 0.62 0.28 0.62 0.28 0.775 0.09 0.775 0.09 0.275 0.16 0.275 0.16 0.115 0.11 0.115 0.11 0.225 0.04 0.225 0.04 0.825 0.11 0.825 0.11 0.95 ;
  END
END BUF_X2P5B_A12TUL_C35

MACRO NAND2B_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN NAND2B_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.23 0.725 0.23 0.55 0.175 0.55 0.175 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.008575 ;
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0238 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.045 0.43 0.875 0.635 0.875 0.635 0.195 0.575 0.195 0.575 0.09 0.505 0.09 0.505 0.27 0.58 0.27 0.58 0.825 0.38 0.825 0.38 1.045 ;
    END
    ANTENNADIFFAREA 0.05775 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.87 0.235 0.87 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.18 1.085 0.18 1.015 0.075 1.015 0.075 0.375 0.445 0.375 0.445 0.69 0.495 0.69 0.495 0.325 0.17 0.325 0.17 0.095 0.1 0.095 0.1 0.325 0.025 0.325 0.025 1.085 ;
  END
END NAND2B_X1M_A12TUL_C35

MACRO CGENI_X1M_A12TH_C35
  CLASS CORE ;
  FOREIGN CGENI_X1M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.495 0.58 0.495 0.58 0.625 0.24 0.625 0.24 0.525 0.16 0.525 0.16 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.575 0.53 0.505 0.365 0.505 0.365 0.425 0.145 0.425 0.145 0.475 0.295 0.475 0.295 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.775 0.77 0.495 0.715 0.495 0.715 0.725 0.55 0.725 0.55 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03045 ;
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 1.005 0.71 0.875 0.905 0.875 0.905 0.325 0.71 0.325 0.71 0.195 0.64 0.195 0.64 0.375 0.85 0.375 0.85 0.825 0.64 0.825 0.64 1.005 ;
    END
    ANTENNADIFFAREA 0.087 ;
  END CON
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.835 0.1 0.835 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.365 0.17 0.035 0.37 0.035 0.37 0.255 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.365 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.845 1.115 0.845 0.93 0.775 0.93 0.775 1.065 0.565 1.065 0.565 0.825 0.245 0.825 0.245 1.015 0.295 1.015 0.295 0.875 0.515 0.875 0.515 1.115 ;
      POLYGON 0.565 0.375 0.565 0.135 0.775 0.135 0.775 0.27 0.845 0.27 0.845 0.085 0.515 0.085 0.515 0.325 0.295 0.325 0.295 0.185 0.245 0.185 0.245 0.375 ;
  END
END CGENI_X1M_A12TH_C35

MACRO BUFH_X2P5M_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUFH_X2P5M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.395 0.475 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0322 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 0.77 0.875 0.77 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.185 0.38 0.185 0.38 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.133875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 0.945 0.505 0.945 0.505 1.165 0.305 1.165 0.305 0.925 0.235 0.925 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.355 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.355 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 0.98 0.16 0.855 0.33 0.855 0.33 0.59 0.56 0.59 0.56 0.61 0.65 0.61 0.65 0.54 0.28 0.54 0.28 0.805 0.09 0.805 0.09 0.355 0.16 0.355 0.16 0.165 0.11 0.165 0.11 0.305 0.04 0.305 0.04 0.855 0.11 0.855 0.11 0.98 ;
  END
END BUFH_X2P5M_A12TUL_C35

MACRO NOR2_X0P5A_A12TL_C35
  CLASS CORE ;
  FOREIGN NOR2_X0P5A_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.54 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.365 0.425 0.145 0.425 0.145 0.475 0.31 0.475 0.31 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.44 1.105 0.44 1.005 0.5 1.005 0.5 0.225 0.295 0.225 0.295 0.145 0.245 0.145 0.245 0.275 0.445 0.275 0.445 0.925 0.37 0.925 0.37 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
      LAYER M1 ;
        POLYGON 0.54 1.235 0.54 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.54 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.205 0.17 0.035 0.365 0.035 0.365 0.17 0.445 0.17 0.445 0.035 0.54 0.035 0.54 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.205 ;
      LAYER M2 ;
        RECT 0 -0.065 0.54 0.065 ;
    END
  END VSS
END NOR2_X0P5A_A12TL_C35

MACRO OA21A1OI2_X4M_A12TUL_C35
  CLASS CORE ;
  FOREIGN OA21A1OI2_X4M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.43 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.175 0.705 1.175 0.425 0.715 0.425 0.715 0.555 0.635 0.555 0.635 0.425 0.175 0.425 0.175 0.705 0.23 0.705 0.23 0.475 0.58 0.475 0.58 0.605 0.77 0.605 0.77 0.475 1.12 0.475 1.12 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.905 0.775 0.905 0.605 1.07 0.605 1.07 0.525 0.83 0.525 0.83 0.725 0.515 0.725 0.515 0.525 0.28 0.525 0.28 0.605 0.445 0.605 0.445 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.445 0.675 1.445 0.625 1.275 0.625 1.275 0.575 1.745 0.575 1.745 0.425 1.63 0.425 1.63 0.475 1.695 0.475 1.695 0.525 1.225 0.525 1.225 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1288 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 2.12 0.675 2.12 0.575 2.285 0.575 2.285 0.425 2.17 0.425 2.17 0.475 2.235 0.475 2.235 0.525 1.86 0.525 1.86 0.485 1.795 0.485 1.795 0.575 2.07 0.575 2.07 0.625 1.9 0.625 1.9 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.102375 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.925 1.005 1.925 0.875 2.135 0.875 2.135 1 2.185 1 2.185 0.875 2.39 0.875 2.39 0.325 2.185 0.325 2.185 0.18 2.135 0.18 2.135 0.325 1.915 0.325 1.915 0.17 1.865 0.17 1.865 0.325 1.645 0.325 1.645 0.2 1.595 0.2 1.595 0.325 1.385 0.325 1.385 0.195 1.315 0.195 1.315 0.375 2.335 0.375 2.335 0.825 1.855 0.825 1.855 1.005 ;
    END
    ANTENNADIFFAREA 0.235625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
        RECT 2.135 1.175 2.185 1.225 ;
        RECT 2.27 1.175 2.32 1.225 ;
      LAYER M1 ;
        POLYGON 2.43 1.235 2.43 1.165 1.655 1.165 1.655 0.945 1.585 0.945 1.585 1.165 1.385 1.165 1.385 0.945 1.315 0.945 1.315 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.43 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
        RECT 2.135 -0.025 2.185 0.025 ;
        RECT 2.27 -0.025 2.32 0.025 ;
      LAYER M1 ;
        POLYGON 2.33 0.27 2.33 0.035 2.43 0.035 2.43 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.505 0.035 0.505 0.255 0.575 0.255 0.575 0.035 0.775 0.035 0.775 0.255 0.845 0.255 0.845 0.035 1.045 0.035 1.045 0.255 1.115 0.255 1.115 0.035 1.99 0.035 1.99 0.255 2.06 0.255 2.06 0.035 2.26 0.035 2.26 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 2.43 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 2.33 1.115 2.33 0.93 2.26 0.93 2.26 1.065 2.05 1.065 2.05 0.94 2 0.94 2 1.065 1.78 1.065 1.78 0.825 0.11 0.825 0.11 1.015 0.16 1.015 0.16 0.875 0.65 0.875 0.65 1 0.7 1 0.7 0.875 1.19 0.875 1.19 1 1.24 1 1.24 0.875 1.46 0.875 1.46 1 1.51 1 1.51 0.875 1.73 0.875 1.73 1.115 ;
      POLYGON 1.24 0.375 1.24 0.135 1.46 0.135 1.46 0.26 1.51 0.26 1.51 0.135 1.72 0.135 1.72 0.27 1.79 0.27 1.79 0.085 1.19 0.085 1.19 0.325 0.97 0.325 0.97 0.2 0.92 0.2 0.92 0.325 0.7 0.325 0.7 0.2 0.65 0.2 0.65 0.325 0.43 0.325 0.43 0.2 0.38 0.2 0.38 0.325 0.16 0.325 0.16 0.185 0.11 0.185 0.11 0.375 ;
  END
END OA21A1OI2_X4M_A12TUL_C35

MACRO NAND4BB_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN NAND4BB_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.945 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.725 0.235 0.575 0.365 0.575 0.365 0.525 0.145 0.525 0.145 0.575 0.165 0.575 0.165 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.665 0.31 0.665 0.31 0.805 0.15 0.805 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END BN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.675 0.645 0.425 0.415 0.425 0.415 0.475 0.565 0.475 0.565 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.565 0.435 0.565 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.835 1.095 0.835 0.975 0.905 0.975 0.905 0.195 0.845 0.195 0.845 0.09 0.775 0.09 0.775 0.27 0.85 0.27 0.85 0.925 0.515 0.925 0.515 1.085 0.565 1.085 0.565 0.975 0.785 0.975 0.785 1.095 ;
    END
    ANTENNADIFFAREA 0.041125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
      LAYER M1 ;
        POLYGON 0.945 1.235 0.945 1.165 0.71 1.165 0.71 1.035 0.64 1.035 0.64 1.165 0.44 1.165 0.44 0.94 0.37 0.94 0.37 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.945 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.255 0.44 0.035 0.945 0.035 0.945 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.945 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.17 1.11 0.17 0.93 0.075 0.93 0.075 0.375 0.715 0.375 0.715 0.515 0.77 0.515 0.77 0.325 0.305 0.325 0.305 0.09 0.235 0.09 0.235 0.325 0.025 0.325 0.025 0.98 0.1 0.98 0.1 1.11 ;
  END
END NAND4BB_X0P5M_A12TUH_C35

MACRO XNOR2_X0P7M_A12TUL_C35
  CLASS CORE ;
  FOREIGN XNOR2_X0P7M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.08 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.19 0.725 0.24 0.775 ;
        RECT 0.475 0.725 0.605 0.775 ;
      LAYER M1 ;
        POLYGON 0.65 0.775 0.65 0.53 0.57 0.53 0.57 0.725 0.43 0.725 0.43 0.775 ;
        RECT 0.18 0.505 0.25 0.825 ;
      LAYER M2 ;
        RECT 0.14 0.725 0.655 0.775 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0065 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02555 LAYER M1 ;
    ANTENNAGATEAREA 0.0546 LAYER M2 ;
    ANTENNAGATEAREA 0.0546 LAYER M3 ;
    ANTENNAGATEAREA 0.0546 LAYER M4 ;
    ANTENNAGATEAREA 0.0546 LAYER M5 ;
    ANTENNAGATEAREA 0.0546 LAYER M6 ;
    ANTENNAGATEAREA 0.0546 LAYER M7 ;
    ANTENNAGATEAREA 0.0546 LAYER M8 ;
    ANTENNAGATEAREA 0.0546 LAYER AP ;
    ANTENNAMAXAREACAR 1.041096 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.2544033 LAYER VIA1 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.935 0.675 0.935 0.605 0.905 0.605 0.905 0.465 0.85 0.465 0.85 0.605 0.715 0.605 0.715 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0308 ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.005 0.575 0.875 1.04 0.875 1.04 0.325 0.72 0.325 0.72 0.3 0.63 0.3 0.63 0.375 0.985 0.375 0.985 0.825 0.505 0.825 0.505 1.005 ;
    END
    ANTENNADIFFAREA 0.079 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
      LAYER M1 ;
        POLYGON 1.08 1.235 1.08 1.165 0.98 1.165 0.98 0.93 0.91 0.93 0.91 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.08 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
      LAYER M1 ;
        POLYGON 0.98 0.27 0.98 0.035 1.08 0.035 1.08 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 0.91 0.035 0.91 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.08 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.845 1.11 0.845 0.93 0.775 0.93 0.775 1.06 0.71 1.06 0.71 0.93 0.64 0.93 0.64 1.06 0.43 1.06 0.43 0.825 0.36 0.825 0.36 0.375 0.565 0.375 0.565 0.25 0.85 0.25 0.85 0.09 0.77 0.09 0.77 0.2 0.515 0.2 0.515 0.325 0.31 0.325 0.31 0.875 0.38 0.875 0.38 1.11 ;
      POLYGON 0.16 1.085 0.16 0.895 0.13 0.895 0.13 0.41 0.16 0.41 0.16 0.22 0.11 0.22 0.11 0.36 0.08 0.36 0.08 0.95 0.11 0.95 0.11 1.085 ;
      POLYGON 0.5 0.6 0.5 0.475 0.71 0.475 0.71 0.54 0.78 0.54 0.78 0.425 0.435 0.425 0.435 0.6 ;
      POLYGON 0.44 0.27 0.44 0.15 0.595 0.15 0.595 0.09 0.37 0.09 0.37 0.27 ;
    LAYER M2 ;
      RECT 0.04 0.425 0.665 0.475 ;
    LAYER VIA1 ;
      RECT 0.485 0.425 0.615 0.475 ;
      RECT 0.08 0.425 0.13 0.475 ;
  END
END XNOR2_X0P7M_A12TUL_C35

MACRO BUF_X1P4B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X1P4B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.495 0.395 0.495 0.395 0.425 0.175 0.425 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01505 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.015 0.43 0.875 0.635 0.875 0.635 0.225 0.43 0.225 0.43 0.12 0.38 0.12 0.38 0.275 0.58 0.275 0.58 0.825 0.38 0.825 0.38 1.015 ;
    END
    ANTENNADIFFAREA 0.051 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.575 1.165 0.575 0.93 0.505 0.93 0.505 1.165 0.305 1.165 0.305 0.895 0.235 0.895 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.195 0.305 0.035 0.5 0.035 0.5 0.17 0.58 0.17 0.58 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.195 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.02 0.16 0.825 0.33 0.825 0.33 0.735 0.495 0.735 0.495 0.545 0.445 0.545 0.445 0.685 0.28 0.685 0.28 0.775 0.09 0.775 0.09 0.18 0.175 0.18 0.175 0.1 0.04 0.1 0.04 0.825 0.11 0.825 0.11 1.02 ;
  END
END BUF_X1P4B_A12TUL_C35

MACRO NAND4_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN NAND4_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.495 0.435 0.495 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.595 0.31 0.595 0.31 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.175 0.475 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.58 1.115 0.58 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.23 0.925 0.23 1.115 0.31 1.115 0.31 0.975 0.5 0.975 0.5 1.115 ;
    END
    ANTENNADIFFAREA 0.03725 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 1.04 0.37 1.04 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.29 0.17 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.29 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND4_X0P5M_A12TUH_C35

MACRO CGENCON_X1M_A12TUL_C35
  CLASS CORE ;
  FOREIGN CGENCON_X1M_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 2.16 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.53 0.495 0.53 0.425 0.305 0.425 0.305 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0287 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.725 0.525 0.775 0.575 ;
        RECT 0.98 0.525 1.03 0.575 ;
        RECT 1.245 0.525 1.295 0.575 ;
      LAYER M1 ;
        POLYGON 0.785 0.7 0.785 0.595 0.795 0.595 0.795 0.505 0.705 0.505 0.705 0.7 ;
        POLYGON 1.05 0.7 1.05 0.505 0.96 0.505 0.96 0.595 0.97 0.595 0.97 0.7 ;
        RECT 1.235 0.445 1.305 0.755 ;
      LAYER M2 ;
        RECT 0.675 0.525 1.345 0.575 ;
    END
    ANTENNAPARTIALMETALAREA 0 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 0 LAYER M8 ;
    ANTENNAPARTIALMETALAREA 0 LAYER AP ;
    ANTENNAPARTIALCUTAREA 0.0025 LAYER VIA1 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015575 LAYER M1 ;
    ANTENNAGATEAREA 0.0616 LAYER M2 ;
    ANTENNAGATEAREA 0.0616 LAYER M3 ;
    ANTENNAGATEAREA 0.0616 LAYER M4 ;
    ANTENNAGATEAREA 0.0616 LAYER M5 ;
    ANTENNAGATEAREA 0.0616 LAYER M6 ;
    ANTENNAGATEAREA 0.0616 LAYER M7 ;
    ANTENNAGATEAREA 0.0616 LAYER M8 ;
    ANTENNAGATEAREA 0.0616 LAYER AP ;
    ANTENNAMAXAREACAR 1.05939 LAYER M2 ;
    ANTENNAMAXAREACAR 0 LAYER M3 ;
    ANTENNAMAXAREACAR 0 LAYER M4 ;
    ANTENNAMAXAREACAR 0 LAYER M5 ;
    ANTENNAMAXAREACAR 0 LAYER M6 ;
    ANTENNAMAXAREACAR 0 LAYER M7 ;
    ANTENNAMAXAREACAR 0 LAYER M8 ;
    ANTENNAMAXAREACAR 0 LAYER AP ;
    ANTENNAMAXCUTCAR 0.1605138 LAYER VIA1 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.92 0.495 1.99 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.028 ;
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 1.645 1.015 1.645 0.875 1.85 0.875 1.85 0.425 1.675 0.425 1.675 0.41 1.525 0.41 1.525 0.475 1.795 0.475 1.795 0.825 1.595 0.825 1.595 1.015 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END CON
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
        RECT 1.19 1.175 1.24 1.225 ;
        RECT 1.325 1.175 1.375 1.225 ;
        RECT 1.46 1.175 1.51 1.225 ;
        RECT 1.595 1.175 1.645 1.225 ;
        RECT 1.73 1.175 1.78 1.225 ;
        RECT 1.865 1.175 1.915 1.225 ;
        RECT 2 1.175 2.05 1.225 ;
      LAYER M1 ;
        POLYGON 2.16 1.235 2.16 1.165 2.065 1.165 2.065 1.03 1.985 1.03 1.985 1.165 1.25 1.165 1.25 0.89 1.18 0.89 1.18 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 2.16 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
        RECT 1.19 -0.025 1.24 0.025 ;
        RECT 1.325 -0.025 1.375 0.025 ;
        RECT 1.46 -0.025 1.51 0.025 ;
        RECT 1.595 -0.025 1.645 0.025 ;
        RECT 1.73 -0.025 1.78 0.025 ;
        RECT 1.865 -0.025 1.915 0.025 ;
        RECT 2 -0.025 2.05 0.025 ;
      LAYER M1 ;
        POLYGON 2.06 0.27 2.06 0.035 2.16 0.035 2.16 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 0.305 0.255 0.305 0.035 1.31 0.035 1.31 0.26 1.39 0.26 1.39 0.035 1.99 0.035 1.99 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 2.16 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 1.79 1.105 1.79 0.975 1.865 0.975 1.865 1.1 1.915 1.1 1.915 0.975 2.12 0.975 2.12 0.325 1.915 0.325 1.915 0.085 1.445 0.085 1.445 0.26 1.525 0.26 1.525 0.135 1.865 0.135 1.865 0.375 2.07 0.375 2.07 0.925 1.72 0.925 1.72 1.105 ;
      POLYGON 1.105 1.045 1.105 0.82 1.17 0.82 1.17 0.41 1.135 0.41 1.135 0.305 0.865 0.305 0.865 0.285 0.755 0.285 0.755 0.355 1.085 0.355 1.085 0.46 1.12 0.46 1.12 0.77 1.055 0.77 1.055 0.995 0.63 0.995 0.63 0.955 0.43 0.955 0.43 0.835 0.095 0.835 0.095 0.27 0.17 0.27 0.17 0.09 0.1 0.09 0.1 0.22 0.045 0.22 0.045 0.885 0.11 0.885 0.11 1.01 0.16 1.01 0.16 0.885 0.38 0.885 0.38 1.005 0.58 1.005 0.58 1.045 ;
      POLYGON 1.51 1.025 1.51 0.835 1.415 0.835 1.415 0.36 1.795 0.36 1.795 0.2 1.715 0.2 1.715 0.31 1.24 0.31 1.24 0.085 0.555 0.085 0.555 0.135 1.19 0.135 1.19 0.36 1.365 0.36 1.365 0.835 1.325 0.835 1.325 1.025 1.375 1.025 1.375 0.885 1.46 0.885 1.46 1.025 ;
      POLYGON 0.98 0.935 0.98 0.755 0.9 0.755 0.9 0.455 1 0.455 1 0.405 0.85 0.405 0.85 0.805 0.91 0.805 0.91 0.935 ;
      POLYGON 0.85 0.935 0.85 0.855 0.54 0.855 0.54 0.735 0.225 0.735 0.225 0.375 0.46 0.375 0.46 0.355 0.61 0.355 0.61 0.235 1.035 0.235 1.035 0.255 1.125 0.255 1.125 0.185 0.56 0.185 0.56 0.305 0.43 0.305 0.43 0.2 0.38 0.2 0.38 0.325 0.175 0.325 0.175 0.785 0.49 0.785 0.49 0.905 0.77 0.905 0.77 0.935 ;
      POLYGON 0.73 0.805 0.73 0.755 0.645 0.755 0.645 0.455 0.73 0.455 0.73 0.405 0.595 0.405 0.595 0.625 0.435 0.625 0.435 0.675 0.595 0.675 0.595 0.805 ;
      POLYGON 1.59 0.775 1.59 0.525 1.51 0.525 1.51 0.705 1.47 0.705 1.47 0.775 ;
      RECT 1.65 0.525 1.73 0.765 ;
    LAYER M2 ;
      RECT 0.8 0.725 1.605 0.775 ;
      RECT 0.425 0.625 1.765 0.675 ;
    LAYER VIA1 ;
      RECT 1.505 0.725 1.555 0.775 ;
      RECT 0.85 0.725 0.9 0.775 ;
      RECT 1.665 0.625 1.715 0.675 ;
      RECT 0.475 0.625 0.605 0.675 ;
  END
END CGENCON_X1M_A12TUL_C35

MACRO NAND4_X0P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN NAND4_X0P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.775 0.635 0.725 0.505 0.725 0.505 0.495 0.435 0.495 0.435 0.705 0.415 0.705 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.875 0.395 0.825 0.365 0.825 0.365 0.595 0.31 0.595 0.31 0.825 0.15 0.825 0.15 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.23 0.705 0.23 0.475 0.365 0.475 0.365 0.425 0.145 0.425 0.145 0.475 0.175 0.475 0.175 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01155 ;
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.58 1.115 0.58 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.23 0.925 0.23 1.115 0.31 1.115 0.31 0.975 0.5 0.975 0.5 1.115 ;
    END
    ANTENNADIFFAREA 0.03725 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.715 1.165 0.715 1.03 0.635 1.03 0.635 1.165 0.44 1.165 0.44 1.04 0.37 1.04 0.37 1.165 0.17 1.165 0.17 1.03 0.1 1.03 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.29 0.17 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.29 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
END NAND4_X0P5M_A12TH_C35

MACRO BUF_X5B_A12TUL_C35
  CLASS CORE ;
  FOREIGN BUF_X5B_A12TUL_C35 ;
  ORIGIN 0 0 ;
  SIZE 1.215 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.575 0.395 0.425 0.145 0.425 0.145 0.475 0.345 0.475 0.345 0.525 0.145 0.525 0.145 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03605 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.015 0.565 0.875 0.785 0.875 0.785 1 0.835 1 0.835 0.875 1.055 0.875 1.055 1 1.105 1 1.105 0.875 1.175 0.875 1.175 0.325 1.115 0.325 1.115 0.09 1.045 0.09 1.045 0.325 0.835 0.325 0.835 0.095 0.785 0.095 0.785 0.325 0.565 0.325 0.565 0.095 0.515 0.095 0.515 0.375 1.12 0.375 1.12 0.825 0.515 0.825 0.515 1.015 ;
    END
    ANTENNADIFFAREA 0.198 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
        RECT 0.785 1.175 0.835 1.225 ;
        RECT 0.92 1.175 0.97 1.225 ;
        RECT 1.055 1.175 1.105 1.225 ;
      LAYER M1 ;
        POLYGON 1.215 1.235 1.215 1.165 0.98 1.165 0.98 0.945 0.91 0.945 0.91 1.165 0.71 1.165 0.71 0.945 0.64 0.945 0.64 1.165 0.44 1.165 0.44 0.845 0.37 0.845 0.37 1.165 0.17 1.165 0.17 0.845 0.1 0.845 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 1.215 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
        RECT 0.785 -0.025 0.835 0.025 ;
        RECT 0.92 -0.025 0.97 0.025 ;
        RECT 1.055 -0.025 1.105 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.27 0.44 0.035 0.64 0.035 0.64 0.255 0.71 0.255 0.71 0.035 0.91 0.035 0.91 0.255 0.98 0.255 0.98 0.035 1.215 0.035 1.215 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.195 0.17 0.195 0.17 0.035 0.37 0.035 0.37 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 1.215 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.295 0.95 0.295 0.775 0.495 0.775 0.495 0.555 0.965 0.555 0.965 0.575 1.055 0.575 1.055 0.505 0.445 0.505 0.445 0.725 0.075 0.725 0.075 0.325 0.295 0.325 0.295 0.12 0.245 0.12 0.245 0.275 0.025 0.275 0.025 0.775 0.245 0.775 0.245 0.95 ;
  END
END BUF_X5B_A12TUL_C35

MACRO AO21A1AI2_X0P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN AO21A1AI2_X0P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.775 0.365 0.725 0.24 0.725 0.24 0.525 0.16 0.525 0.16 0.725 0.145 0.725 0.145 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.495 0.395 0.495 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.635 0.675 0.635 0.625 0.5 0.625 0.5 0.465 0.445 0.465 0.445 0.605 0.415 0.605 0.415 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.016275 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.575 0.645 0.325 0.415 0.325 0.415 0.375 0.565 0.375 0.565 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012775 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 1.07 0.565 0.875 0.77 0.875 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.275 0.715 0.275 0.715 0.825 0.515 0.825 0.515 1.07 ;
    END
    ANTENNADIFFAREA 0.03875 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 1.005 0.64 1.005 0.64 1.165 0.305 1.165 0.305 0.945 0.235 0.945 0.235 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.44 0.165 0.44 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.37 0.035 0.37 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.16 1.07 0.16 0.875 0.38 0.875 0.38 1.06 0.43 1.06 0.43 0.825 0.11 0.825 0.11 1.07 ;
      POLYGON 0.575 0.275 0.575 0.095 0.505 0.095 0.505 0.225 0.17 0.225 0.17 0.09 0.1 0.09 0.1 0.275 ;
  END
END AO21A1AI2_X0P5M_A12TH_C35

MACRO OAI22_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN OAI22_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.44 0.495 0.44 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.775 0.64 0.565 0.57 0.565 0.57 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.015225 ;
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.43 1.06 0.43 0.875 0.77 0.875 0.77 0.325 0.58 0.325 0.58 0.185 0.5 0.185 0.5 0.375 0.715 0.375 0.715 0.825 0.38 0.825 0.38 1.06 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.71 1.165 0.71 0.925 0.64 0.925 0.64 1.165 0.17 1.165 0.17 0.885 0.1 0.885 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.165 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.165 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.44 0.275 0.44 0.135 0.65 0.135 0.65 0.22 0.7 0.22 0.7 0.085 0.37 0.085 0.37 0.225 0.16 0.225 0.16 0.11 0.11 0.11 0.11 0.275 ;
  END
END OAI22_X0P5M_A12TL_C35

MACRO AOI31_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN AOI31_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.635 0.5 0.475 0.635 0.475 0.635 0.425 0.415 0.425 0.415 0.495 0.445 0.495 0.445 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.395 0.675 0.395 0.605 0.365 0.605 0.365 0.465 0.31 0.465 0.31 0.625 0.15 0.625 0.15 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.575 0.24 0.375 0.365 0.375 0.365 0.325 0.145 0.325 0.145 0.375 0.16 0.375 0.16 0.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.645 0.775 0.645 0.525 0.565 0.525 0.565 0.725 0.415 0.725 0.415 0.775 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.013125 ;
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 1.065 0.7 0.905 0.77 0.905 0.77 0.325 0.575 0.325 0.575 0.09 0.505 0.09 0.505 0.27 0.525 0.27 0.525 0.375 0.715 0.375 0.715 0.855 0.65 0.855 0.65 1.065 ;
    END
    ANTENNADIFFAREA 0.038125 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.44 1.165 0.44 0.945 0.37 0.945 0.37 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.64 0.035 0.64 0.175 0.71 0.175 0.71 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.565 1.055 0.565 0.825 0.245 0.825 0.245 1.055 0.295 1.055 0.295 0.875 0.515 0.875 0.515 1.055 ;
  END
END AOI31_X0P5M_A12TL_C35

MACRO NOR3_X0P5M_A12TUH_C35
  CLASS CORE ;
  FOREIGN NOR3_X0P5M_A12TUH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.875 0.5 0.595 0.445 0.595 0.445 0.825 0.28 0.825 0.28 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.225 0.58 0.225 0.58 0.085 0.5 0.085 0.5 0.225 0.305 0.225 0.305 0.095 0.235 0.095 0.235 0.275 0.58 0.275 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END NOR3_X0P5M_A12TUH_C35

MACRO OAI211_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN OAI211_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.81 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.635 0.365 0.475 0.395 0.475 0.395 0.425 0.15 0.425 0.15 0.475 0.31 0.475 0.31 0.635 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.875 0.365 0.825 0.23 0.825 0.23 0.595 0.175 0.595 0.175 0.825 0.145 0.825 0.145 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0154 ;
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.64 0.595 0.64 0.395 0.58 0.395 0.58 0.525 0.415 0.525 0.415 0.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.875 0.665 0.705 0.415 0.705 0.415 0.775 0.615 0.775 0.615 0.825 0.55 0.825 0.55 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.011025 ;
  END C0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 1.11 0.715 0.975 0.77 0.975 0.77 0.195 0.71 0.195 0.71 0.09 0.64 0.09 0.64 0.27 0.715 0.27 0.715 0.925 0.37 0.925 0.37 1.105 0.44 1.105 0.44 0.975 0.635 0.975 0.635 1.11 ;
    END
    ANTENNADIFFAREA 0.0435 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
        RECT 0.65 1.175 0.7 1.225 ;
      LAYER M1 ;
        POLYGON 0.81 1.235 0.81 1.165 0.575 1.165 0.575 1.04 0.505 1.04 0.505 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.81 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
        RECT 0.65 -0.025 0.7 0.025 ;
      LAYER M1 ;
        POLYGON 0.305 0.255 0.305 0.035 0.81 0.035 0.81 -0.035 0 -0.035 0 0.035 0.235 0.035 0.235 0.255 ;
      LAYER M2 ;
        RECT 0 -0.065 0.81 0.065 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      POLYGON 0.43 0.375 0.43 0.095 0.38 0.095 0.38 0.325 0.17 0.325 0.17 0.09 0.1 0.09 0.1 0.27 0.12 0.27 0.12 0.375 ;
  END
END OAI211_X0P5M_A12TL_C35

MACRO INV_X0P5M_A12TL_C35
  CLASS CORE ;
  FOREIGN INV_X0P5M_A12TL_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.405 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.175 0.395 0.23 0.805 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.01645 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 1.065 0.295 0.925 0.365 0.925 0.365 0.195 0.305 0.195 0.305 0.09 0.235 0.09 0.235 0.27 0.31 0.27 0.31 0.875 0.245 0.875 0.245 1.065 ;
    END
    ANTENNADIFFAREA 0.03525 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
      LAYER M1 ;
        POLYGON 0.405 1.235 0.405 1.165 0.17 1.165 0.17 0.88 0.1 0.88 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.405 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.27 0.17 0.035 0.405 0.035 0.405 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.27 ;
      LAYER M2 ;
        RECT 0 -0.065 0.405 0.065 ;
    END
  END VSS
END INV_X0P5M_A12TL_C35

MACRO NOR3_X0P5M_A12TH_C35
  CLASS CORE ;
  FOREIGN NOR3_X0P5M_A12TH_C35 ;
  ORIGIN 0 0 ;
  SIZE 0.675 BY 1.2 ;
  SYMMETRY X Y ;
  SITE sc12mc_cln28hpm ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.875 0.5 0.595 0.445 0.595 0.445 0.825 0.28 0.825 0.28 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.535 0.365 0.375 0.395 0.375 0.395 0.325 0.15 0.325 0.15 0.375 0.305 0.375 0.305 0.535 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.675 0.365 0.625 0.235 0.625 0.235 0.465 0.165 0.465 0.165 0.625 0.145 0.625 0.145 0.675 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.012425 ;
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        POLYGON 0.575 1.105 0.575 1.005 0.635 1.005 0.635 0.225 0.58 0.225 0.58 0.085 0.5 0.085 0.5 0.225 0.305 0.225 0.305 0.095 0.235 0.095 0.235 0.275 0.58 0.275 0.58 0.925 0.505 0.925 0.505 1.105 ;
    END
    ANTENNADIFFAREA 0.036625 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 1.175 0.16 1.225 ;
        RECT 0.245 1.175 0.295 1.225 ;
        RECT 0.38 1.175 0.43 1.225 ;
        RECT 0.515 1.175 0.565 1.225 ;
      LAYER M1 ;
        POLYGON 0.675 1.235 0.675 1.165 0.17 1.165 0.17 0.93 0.1 0.93 0.1 1.165 0 1.165 0 1.235 ;
      LAYER M2 ;
        RECT 0 1.135 0.675 1.265 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER VIA1 ;
        RECT 0.11 -0.025 0.16 0.025 ;
        RECT 0.245 -0.025 0.295 0.025 ;
        RECT 0.38 -0.025 0.43 0.025 ;
        RECT 0.515 -0.025 0.565 0.025 ;
      LAYER M1 ;
        POLYGON 0.17 0.17 0.17 0.035 0.37 0.035 0.37 0.165 0.44 0.165 0.44 0.035 0.675 0.035 0.675 -0.035 0 -0.035 0 0.035 0.1 0.035 0.1 0.17 ;
      LAYER M2 ;
        RECT 0 -0.065 0.675 0.065 ;
    END
  END VSS
END NOR3_X0P5M_A12TH_C35

END LIBRARY
